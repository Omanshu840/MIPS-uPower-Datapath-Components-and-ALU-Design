$date
	Sun May 31 02:15:07 2020
$end
$version
	Icarus Verilog
$end
$timescale
	1s
$end
$scope module tb_uPOWER_ALU_ALUCU $end
$var wire 4 ! ALUControl [3:0] $end
$var wire 1 " Overflow $end
$var wire 64 # Result [63:0] $end
$var wire 1 $ Zero $end
$var reg 2 % ALUOp [1:0] $end
$var reg 6 & OpCode [5:0] $end
$var reg 9 ' XO [8:0] $end
$var reg 64 ( a [63:0] $end
$var reg 64 ) b [63:0] $end
$scope module C $end
$var wire 4 * ALUControl [3:0] $end
$var wire 17 + ALUControlIn [16:0] $end
$var wire 2 , ALUOp [1:0] $end
$var wire 6 - OpCode [5:0] $end
$var wire 9 . XO [8:0] $end
$var reg 4 / ALUCtrl [3:0] $end
$upscope $end
$scope module A $end
$var wire 4 0 ALUOperatn [3:0] $end
$var wire 64 1 CarryOut [63:0] $end
$var wire 1 " Overflow $end
$var wire 64 2 Result [63:0] $end
$var wire 1 3 Set $end
$var wire 1 $ Zero $end
$var wire 64 4 a [63:0] $end
$var wire 64 5 b [63:0] $end
$scope module A0 $end
$var wire 1 6 Ainvert $end
$var wire 1 7 Binvert $end
$var wire 1 8 CarryIn $end
$var wire 1 9 CarryOut $end
$var wire 1 3 Less $end
$var wire 2 : Operation [1:0] $end
$var wire 1 ; Result $end
$var wire 1 < a $end
$var wire 1 = b $end
$var wire 2 > mux0inputs [1:0] $end
$var wire 2 ? mux1inputs [1:0] $end
$var wire 4 @ mux2inputs [3:0] $end
$var wire 1 A w1 $end
$var wire 1 B w2 $end
$scope module P0 $end
$var wire 2 C inputLines [1:0] $end
$var wire 1 A outputLine $end
$var wire 1 6 selectLine $end
$var wire 1 D w1 $end
$var wire 1 E w2 $end
$var wire 1 F w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 G inputLines [1:0] $end
$var wire 1 B outputLine $end
$var wire 1 7 selectLine $end
$var wire 1 H w1 $end
$var wire 1 I w2 $end
$var wire 1 J w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 A a $end
$var wire 1 B b $end
$var wire 1 8 cin $end
$var wire 1 9 cout $end
$var wire 1 K sum $end
$var wire 1 L w1 $end
$var wire 1 M w2 $end
$var wire 1 N w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 O inputLines [3:0] $end
$var wire 1 ; outputLine $end
$var wire 2 P selectLines [1:0] $end
$var wire 2 Q w [1:0] $end
$scope module M0 $end
$var wire 2 R inputLines [1:0] $end
$var wire 1 S outputLine $end
$var wire 1 T selectLine $end
$var wire 1 U w1 $end
$var wire 1 V w2 $end
$var wire 1 W w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 X inputLines [1:0] $end
$var wire 1 Y outputLine $end
$var wire 1 Z selectLine $end
$var wire 1 [ w1 $end
$var wire 1 \ w2 $end
$var wire 1 ] w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 ^ inputLines [1:0] $end
$var wire 1 ; outputLine $end
$var wire 1 _ selectLine $end
$var wire 1 ` w1 $end
$var wire 1 a w2 $end
$var wire 1 b w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A1 $end
$var wire 1 c Ainvert $end
$var wire 1 d Binvert $end
$var wire 1 e CarryIn $end
$var wire 1 f CarryOut $end
$var wire 1 g Less $end
$var wire 2 h Operation [1:0] $end
$var wire 1 i Result $end
$var wire 1 j a $end
$var wire 1 k b $end
$var wire 2 l mux0inputs [1:0] $end
$var wire 2 m mux1inputs [1:0] $end
$var wire 4 n mux2inputs [3:0] $end
$var wire 1 o w1 $end
$var wire 1 p w2 $end
$scope module P0 $end
$var wire 2 q inputLines [1:0] $end
$var wire 1 o outputLine $end
$var wire 1 c selectLine $end
$var wire 1 r w1 $end
$var wire 1 s w2 $end
$var wire 1 t w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 u inputLines [1:0] $end
$var wire 1 p outputLine $end
$var wire 1 d selectLine $end
$var wire 1 v w1 $end
$var wire 1 w w2 $end
$var wire 1 x w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 o a $end
$var wire 1 p b $end
$var wire 1 e cin $end
$var wire 1 f cout $end
$var wire 1 y sum $end
$var wire 1 z w1 $end
$var wire 1 { w2 $end
$var wire 1 | w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 } inputLines [3:0] $end
$var wire 1 i outputLine $end
$var wire 2 ~ selectLines [1:0] $end
$var wire 2 !" w [1:0] $end
$scope module M0 $end
$var wire 2 "" inputLines [1:0] $end
$var wire 1 #" outputLine $end
$var wire 1 $" selectLine $end
$var wire 1 %" w1 $end
$var wire 1 &" w2 $end
$var wire 1 '" w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 (" inputLines [1:0] $end
$var wire 1 )" outputLine $end
$var wire 1 *" selectLine $end
$var wire 1 +" w1 $end
$var wire 1 ," w2 $end
$var wire 1 -" w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 ." inputLines [1:0] $end
$var wire 1 i outputLine $end
$var wire 1 /" selectLine $end
$var wire 1 0" w1 $end
$var wire 1 1" w2 $end
$var wire 1 2" w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A2 $end
$var wire 1 3" Ainvert $end
$var wire 1 4" Binvert $end
$var wire 1 5" CarryIn $end
$var wire 1 6" CarryOut $end
$var wire 1 7" Less $end
$var wire 2 8" Operation [1:0] $end
$var wire 1 9" Result $end
$var wire 1 :" a $end
$var wire 1 ;" b $end
$var wire 2 <" mux0inputs [1:0] $end
$var wire 2 =" mux1inputs [1:0] $end
$var wire 4 >" mux2inputs [3:0] $end
$var wire 1 ?" w1 $end
$var wire 1 @" w2 $end
$scope module P0 $end
$var wire 2 A" inputLines [1:0] $end
$var wire 1 ?" outputLine $end
$var wire 1 3" selectLine $end
$var wire 1 B" w1 $end
$var wire 1 C" w2 $end
$var wire 1 D" w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 E" inputLines [1:0] $end
$var wire 1 @" outputLine $end
$var wire 1 4" selectLine $end
$var wire 1 F" w1 $end
$var wire 1 G" w2 $end
$var wire 1 H" w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 ?" a $end
$var wire 1 @" b $end
$var wire 1 5" cin $end
$var wire 1 6" cout $end
$var wire 1 I" sum $end
$var wire 1 J" w1 $end
$var wire 1 K" w2 $end
$var wire 1 L" w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 M" inputLines [3:0] $end
$var wire 1 9" outputLine $end
$var wire 2 N" selectLines [1:0] $end
$var wire 2 O" w [1:0] $end
$scope module M0 $end
$var wire 2 P" inputLines [1:0] $end
$var wire 1 Q" outputLine $end
$var wire 1 R" selectLine $end
$var wire 1 S" w1 $end
$var wire 1 T" w2 $end
$var wire 1 U" w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 V" inputLines [1:0] $end
$var wire 1 W" outputLine $end
$var wire 1 X" selectLine $end
$var wire 1 Y" w1 $end
$var wire 1 Z" w2 $end
$var wire 1 [" w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 \" inputLines [1:0] $end
$var wire 1 9" outputLine $end
$var wire 1 ]" selectLine $end
$var wire 1 ^" w1 $end
$var wire 1 _" w2 $end
$var wire 1 `" w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A3 $end
$var wire 1 a" Ainvert $end
$var wire 1 b" Binvert $end
$var wire 1 c" CarryIn $end
$var wire 1 d" CarryOut $end
$var wire 1 e" Less $end
$var wire 2 f" Operation [1:0] $end
$var wire 1 g" Result $end
$var wire 1 h" a $end
$var wire 1 i" b $end
$var wire 2 j" mux0inputs [1:0] $end
$var wire 2 k" mux1inputs [1:0] $end
$var wire 4 l" mux2inputs [3:0] $end
$var wire 1 m" w1 $end
$var wire 1 n" w2 $end
$scope module P0 $end
$var wire 2 o" inputLines [1:0] $end
$var wire 1 m" outputLine $end
$var wire 1 a" selectLine $end
$var wire 1 p" w1 $end
$var wire 1 q" w2 $end
$var wire 1 r" w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 s" inputLines [1:0] $end
$var wire 1 n" outputLine $end
$var wire 1 b" selectLine $end
$var wire 1 t" w1 $end
$var wire 1 u" w2 $end
$var wire 1 v" w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 m" a $end
$var wire 1 n" b $end
$var wire 1 c" cin $end
$var wire 1 d" cout $end
$var wire 1 w" sum $end
$var wire 1 x" w1 $end
$var wire 1 y" w2 $end
$var wire 1 z" w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 {" inputLines [3:0] $end
$var wire 1 g" outputLine $end
$var wire 2 |" selectLines [1:0] $end
$var wire 2 }" w [1:0] $end
$scope module M0 $end
$var wire 2 ~" inputLines [1:0] $end
$var wire 1 !# outputLine $end
$var wire 1 "# selectLine $end
$var wire 1 ## w1 $end
$var wire 1 $# w2 $end
$var wire 1 %# w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 &# inputLines [1:0] $end
$var wire 1 '# outputLine $end
$var wire 1 (# selectLine $end
$var wire 1 )# w1 $end
$var wire 1 *# w2 $end
$var wire 1 +# w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 ,# inputLines [1:0] $end
$var wire 1 g" outputLine $end
$var wire 1 -# selectLine $end
$var wire 1 .# w1 $end
$var wire 1 /# w2 $end
$var wire 1 0# w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A4 $end
$var wire 1 1# Ainvert $end
$var wire 1 2# Binvert $end
$var wire 1 3# CarryIn $end
$var wire 1 4# CarryOut $end
$var wire 1 5# Less $end
$var wire 2 6# Operation [1:0] $end
$var wire 1 7# Result $end
$var wire 1 8# a $end
$var wire 1 9# b $end
$var wire 2 :# mux0inputs [1:0] $end
$var wire 2 ;# mux1inputs [1:0] $end
$var wire 4 <# mux2inputs [3:0] $end
$var wire 1 =# w1 $end
$var wire 1 ># w2 $end
$scope module P0 $end
$var wire 2 ?# inputLines [1:0] $end
$var wire 1 =# outputLine $end
$var wire 1 1# selectLine $end
$var wire 1 @# w1 $end
$var wire 1 A# w2 $end
$var wire 1 B# w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 C# inputLines [1:0] $end
$var wire 1 ># outputLine $end
$var wire 1 2# selectLine $end
$var wire 1 D# w1 $end
$var wire 1 E# w2 $end
$var wire 1 F# w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 =# a $end
$var wire 1 ># b $end
$var wire 1 3# cin $end
$var wire 1 4# cout $end
$var wire 1 G# sum $end
$var wire 1 H# w1 $end
$var wire 1 I# w2 $end
$var wire 1 J# w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 K# inputLines [3:0] $end
$var wire 1 7# outputLine $end
$var wire 2 L# selectLines [1:0] $end
$var wire 2 M# w [1:0] $end
$scope module M0 $end
$var wire 2 N# inputLines [1:0] $end
$var wire 1 O# outputLine $end
$var wire 1 P# selectLine $end
$var wire 1 Q# w1 $end
$var wire 1 R# w2 $end
$var wire 1 S# w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 T# inputLines [1:0] $end
$var wire 1 U# outputLine $end
$var wire 1 V# selectLine $end
$var wire 1 W# w1 $end
$var wire 1 X# w2 $end
$var wire 1 Y# w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 Z# inputLines [1:0] $end
$var wire 1 7# outputLine $end
$var wire 1 [# selectLine $end
$var wire 1 \# w1 $end
$var wire 1 ]# w2 $end
$var wire 1 ^# w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A5 $end
$var wire 1 _# Ainvert $end
$var wire 1 `# Binvert $end
$var wire 1 a# CarryIn $end
$var wire 1 b# CarryOut $end
$var wire 1 c# Less $end
$var wire 2 d# Operation [1:0] $end
$var wire 1 e# Result $end
$var wire 1 f# a $end
$var wire 1 g# b $end
$var wire 2 h# mux0inputs [1:0] $end
$var wire 2 i# mux1inputs [1:0] $end
$var wire 4 j# mux2inputs [3:0] $end
$var wire 1 k# w1 $end
$var wire 1 l# w2 $end
$scope module P0 $end
$var wire 2 m# inputLines [1:0] $end
$var wire 1 k# outputLine $end
$var wire 1 _# selectLine $end
$var wire 1 n# w1 $end
$var wire 1 o# w2 $end
$var wire 1 p# w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 q# inputLines [1:0] $end
$var wire 1 l# outputLine $end
$var wire 1 `# selectLine $end
$var wire 1 r# w1 $end
$var wire 1 s# w2 $end
$var wire 1 t# w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 k# a $end
$var wire 1 l# b $end
$var wire 1 a# cin $end
$var wire 1 b# cout $end
$var wire 1 u# sum $end
$var wire 1 v# w1 $end
$var wire 1 w# w2 $end
$var wire 1 x# w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 y# inputLines [3:0] $end
$var wire 1 e# outputLine $end
$var wire 2 z# selectLines [1:0] $end
$var wire 2 {# w [1:0] $end
$scope module M0 $end
$var wire 2 |# inputLines [1:0] $end
$var wire 1 }# outputLine $end
$var wire 1 ~# selectLine $end
$var wire 1 !$ w1 $end
$var wire 1 "$ w2 $end
$var wire 1 #$ w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 $$ inputLines [1:0] $end
$var wire 1 %$ outputLine $end
$var wire 1 &$ selectLine $end
$var wire 1 '$ w1 $end
$var wire 1 ($ w2 $end
$var wire 1 )$ w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 *$ inputLines [1:0] $end
$var wire 1 e# outputLine $end
$var wire 1 +$ selectLine $end
$var wire 1 ,$ w1 $end
$var wire 1 -$ w2 $end
$var wire 1 .$ w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A6 $end
$var wire 1 /$ Ainvert $end
$var wire 1 0$ Binvert $end
$var wire 1 1$ CarryIn $end
$var wire 1 2$ CarryOut $end
$var wire 1 3$ Less $end
$var wire 2 4$ Operation [1:0] $end
$var wire 1 5$ Result $end
$var wire 1 6$ a $end
$var wire 1 7$ b $end
$var wire 2 8$ mux0inputs [1:0] $end
$var wire 2 9$ mux1inputs [1:0] $end
$var wire 4 :$ mux2inputs [3:0] $end
$var wire 1 ;$ w1 $end
$var wire 1 <$ w2 $end
$scope module P0 $end
$var wire 2 =$ inputLines [1:0] $end
$var wire 1 ;$ outputLine $end
$var wire 1 /$ selectLine $end
$var wire 1 >$ w1 $end
$var wire 1 ?$ w2 $end
$var wire 1 @$ w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 A$ inputLines [1:0] $end
$var wire 1 <$ outputLine $end
$var wire 1 0$ selectLine $end
$var wire 1 B$ w1 $end
$var wire 1 C$ w2 $end
$var wire 1 D$ w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 ;$ a $end
$var wire 1 <$ b $end
$var wire 1 1$ cin $end
$var wire 1 2$ cout $end
$var wire 1 E$ sum $end
$var wire 1 F$ w1 $end
$var wire 1 G$ w2 $end
$var wire 1 H$ w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 I$ inputLines [3:0] $end
$var wire 1 5$ outputLine $end
$var wire 2 J$ selectLines [1:0] $end
$var wire 2 K$ w [1:0] $end
$scope module M0 $end
$var wire 2 L$ inputLines [1:0] $end
$var wire 1 M$ outputLine $end
$var wire 1 N$ selectLine $end
$var wire 1 O$ w1 $end
$var wire 1 P$ w2 $end
$var wire 1 Q$ w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 R$ inputLines [1:0] $end
$var wire 1 S$ outputLine $end
$var wire 1 T$ selectLine $end
$var wire 1 U$ w1 $end
$var wire 1 V$ w2 $end
$var wire 1 W$ w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 X$ inputLines [1:0] $end
$var wire 1 5$ outputLine $end
$var wire 1 Y$ selectLine $end
$var wire 1 Z$ w1 $end
$var wire 1 [$ w2 $end
$var wire 1 \$ w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A7 $end
$var wire 1 ]$ Ainvert $end
$var wire 1 ^$ Binvert $end
$var wire 1 _$ CarryIn $end
$var wire 1 `$ CarryOut $end
$var wire 1 a$ Less $end
$var wire 2 b$ Operation [1:0] $end
$var wire 1 c$ Result $end
$var wire 1 d$ a $end
$var wire 1 e$ b $end
$var wire 2 f$ mux0inputs [1:0] $end
$var wire 2 g$ mux1inputs [1:0] $end
$var wire 4 h$ mux2inputs [3:0] $end
$var wire 1 i$ w1 $end
$var wire 1 j$ w2 $end
$scope module P0 $end
$var wire 2 k$ inputLines [1:0] $end
$var wire 1 i$ outputLine $end
$var wire 1 ]$ selectLine $end
$var wire 1 l$ w1 $end
$var wire 1 m$ w2 $end
$var wire 1 n$ w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 o$ inputLines [1:0] $end
$var wire 1 j$ outputLine $end
$var wire 1 ^$ selectLine $end
$var wire 1 p$ w1 $end
$var wire 1 q$ w2 $end
$var wire 1 r$ w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 i$ a $end
$var wire 1 j$ b $end
$var wire 1 _$ cin $end
$var wire 1 `$ cout $end
$var wire 1 s$ sum $end
$var wire 1 t$ w1 $end
$var wire 1 u$ w2 $end
$var wire 1 v$ w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 w$ inputLines [3:0] $end
$var wire 1 c$ outputLine $end
$var wire 2 x$ selectLines [1:0] $end
$var wire 2 y$ w [1:0] $end
$scope module M0 $end
$var wire 2 z$ inputLines [1:0] $end
$var wire 1 {$ outputLine $end
$var wire 1 |$ selectLine $end
$var wire 1 }$ w1 $end
$var wire 1 ~$ w2 $end
$var wire 1 !% w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 "% inputLines [1:0] $end
$var wire 1 #% outputLine $end
$var wire 1 $% selectLine $end
$var wire 1 %% w1 $end
$var wire 1 &% w2 $end
$var wire 1 '% w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 (% inputLines [1:0] $end
$var wire 1 c$ outputLine $end
$var wire 1 )% selectLine $end
$var wire 1 *% w1 $end
$var wire 1 +% w2 $end
$var wire 1 ,% w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A8 $end
$var wire 1 -% Ainvert $end
$var wire 1 .% Binvert $end
$var wire 1 /% CarryIn $end
$var wire 1 0% CarryOut $end
$var wire 1 1% Less $end
$var wire 2 2% Operation [1:0] $end
$var wire 1 3% Result $end
$var wire 1 4% a $end
$var wire 1 5% b $end
$var wire 2 6% mux0inputs [1:0] $end
$var wire 2 7% mux1inputs [1:0] $end
$var wire 4 8% mux2inputs [3:0] $end
$var wire 1 9% w1 $end
$var wire 1 :% w2 $end
$scope module P0 $end
$var wire 2 ;% inputLines [1:0] $end
$var wire 1 9% outputLine $end
$var wire 1 -% selectLine $end
$var wire 1 <% w1 $end
$var wire 1 =% w2 $end
$var wire 1 >% w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 ?% inputLines [1:0] $end
$var wire 1 :% outputLine $end
$var wire 1 .% selectLine $end
$var wire 1 @% w1 $end
$var wire 1 A% w2 $end
$var wire 1 B% w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 9% a $end
$var wire 1 :% b $end
$var wire 1 /% cin $end
$var wire 1 0% cout $end
$var wire 1 C% sum $end
$var wire 1 D% w1 $end
$var wire 1 E% w2 $end
$var wire 1 F% w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 G% inputLines [3:0] $end
$var wire 1 3% outputLine $end
$var wire 2 H% selectLines [1:0] $end
$var wire 2 I% w [1:0] $end
$scope module M0 $end
$var wire 2 J% inputLines [1:0] $end
$var wire 1 K% outputLine $end
$var wire 1 L% selectLine $end
$var wire 1 M% w1 $end
$var wire 1 N% w2 $end
$var wire 1 O% w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 P% inputLines [1:0] $end
$var wire 1 Q% outputLine $end
$var wire 1 R% selectLine $end
$var wire 1 S% w1 $end
$var wire 1 T% w2 $end
$var wire 1 U% w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 V% inputLines [1:0] $end
$var wire 1 3% outputLine $end
$var wire 1 W% selectLine $end
$var wire 1 X% w1 $end
$var wire 1 Y% w2 $end
$var wire 1 Z% w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A9 $end
$var wire 1 [% Ainvert $end
$var wire 1 \% Binvert $end
$var wire 1 ]% CarryIn $end
$var wire 1 ^% CarryOut $end
$var wire 1 _% Less $end
$var wire 2 `% Operation [1:0] $end
$var wire 1 a% Result $end
$var wire 1 b% a $end
$var wire 1 c% b $end
$var wire 2 d% mux0inputs [1:0] $end
$var wire 2 e% mux1inputs [1:0] $end
$var wire 4 f% mux2inputs [3:0] $end
$var wire 1 g% w1 $end
$var wire 1 h% w2 $end
$scope module P0 $end
$var wire 2 i% inputLines [1:0] $end
$var wire 1 g% outputLine $end
$var wire 1 [% selectLine $end
$var wire 1 j% w1 $end
$var wire 1 k% w2 $end
$var wire 1 l% w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 m% inputLines [1:0] $end
$var wire 1 h% outputLine $end
$var wire 1 \% selectLine $end
$var wire 1 n% w1 $end
$var wire 1 o% w2 $end
$var wire 1 p% w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 g% a $end
$var wire 1 h% b $end
$var wire 1 ]% cin $end
$var wire 1 ^% cout $end
$var wire 1 q% sum $end
$var wire 1 r% w1 $end
$var wire 1 s% w2 $end
$var wire 1 t% w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 u% inputLines [3:0] $end
$var wire 1 a% outputLine $end
$var wire 2 v% selectLines [1:0] $end
$var wire 2 w% w [1:0] $end
$scope module M0 $end
$var wire 2 x% inputLines [1:0] $end
$var wire 1 y% outputLine $end
$var wire 1 z% selectLine $end
$var wire 1 {% w1 $end
$var wire 1 |% w2 $end
$var wire 1 }% w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 ~% inputLines [1:0] $end
$var wire 1 !& outputLine $end
$var wire 1 "& selectLine $end
$var wire 1 #& w1 $end
$var wire 1 $& w2 $end
$var wire 1 %& w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 && inputLines [1:0] $end
$var wire 1 a% outputLine $end
$var wire 1 '& selectLine $end
$var wire 1 (& w1 $end
$var wire 1 )& w2 $end
$var wire 1 *& w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A10 $end
$var wire 1 +& Ainvert $end
$var wire 1 ,& Binvert $end
$var wire 1 -& CarryIn $end
$var wire 1 .& CarryOut $end
$var wire 1 /& Less $end
$var wire 2 0& Operation [1:0] $end
$var wire 1 1& Result $end
$var wire 1 2& a $end
$var wire 1 3& b $end
$var wire 2 4& mux0inputs [1:0] $end
$var wire 2 5& mux1inputs [1:0] $end
$var wire 4 6& mux2inputs [3:0] $end
$var wire 1 7& w1 $end
$var wire 1 8& w2 $end
$scope module P0 $end
$var wire 2 9& inputLines [1:0] $end
$var wire 1 7& outputLine $end
$var wire 1 +& selectLine $end
$var wire 1 :& w1 $end
$var wire 1 ;& w2 $end
$var wire 1 <& w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 =& inputLines [1:0] $end
$var wire 1 8& outputLine $end
$var wire 1 ,& selectLine $end
$var wire 1 >& w1 $end
$var wire 1 ?& w2 $end
$var wire 1 @& w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 7& a $end
$var wire 1 8& b $end
$var wire 1 -& cin $end
$var wire 1 .& cout $end
$var wire 1 A& sum $end
$var wire 1 B& w1 $end
$var wire 1 C& w2 $end
$var wire 1 D& w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 E& inputLines [3:0] $end
$var wire 1 1& outputLine $end
$var wire 2 F& selectLines [1:0] $end
$var wire 2 G& w [1:0] $end
$scope module M0 $end
$var wire 2 H& inputLines [1:0] $end
$var wire 1 I& outputLine $end
$var wire 1 J& selectLine $end
$var wire 1 K& w1 $end
$var wire 1 L& w2 $end
$var wire 1 M& w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 N& inputLines [1:0] $end
$var wire 1 O& outputLine $end
$var wire 1 P& selectLine $end
$var wire 1 Q& w1 $end
$var wire 1 R& w2 $end
$var wire 1 S& w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 T& inputLines [1:0] $end
$var wire 1 1& outputLine $end
$var wire 1 U& selectLine $end
$var wire 1 V& w1 $end
$var wire 1 W& w2 $end
$var wire 1 X& w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A11 $end
$var wire 1 Y& Ainvert $end
$var wire 1 Z& Binvert $end
$var wire 1 [& CarryIn $end
$var wire 1 \& CarryOut $end
$var wire 1 ]& Less $end
$var wire 2 ^& Operation [1:0] $end
$var wire 1 _& Result $end
$var wire 1 `& a $end
$var wire 1 a& b $end
$var wire 2 b& mux0inputs [1:0] $end
$var wire 2 c& mux1inputs [1:0] $end
$var wire 4 d& mux2inputs [3:0] $end
$var wire 1 e& w1 $end
$var wire 1 f& w2 $end
$scope module P0 $end
$var wire 2 g& inputLines [1:0] $end
$var wire 1 e& outputLine $end
$var wire 1 Y& selectLine $end
$var wire 1 h& w1 $end
$var wire 1 i& w2 $end
$var wire 1 j& w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 k& inputLines [1:0] $end
$var wire 1 f& outputLine $end
$var wire 1 Z& selectLine $end
$var wire 1 l& w1 $end
$var wire 1 m& w2 $end
$var wire 1 n& w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 e& a $end
$var wire 1 f& b $end
$var wire 1 [& cin $end
$var wire 1 \& cout $end
$var wire 1 o& sum $end
$var wire 1 p& w1 $end
$var wire 1 q& w2 $end
$var wire 1 r& w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 s& inputLines [3:0] $end
$var wire 1 _& outputLine $end
$var wire 2 t& selectLines [1:0] $end
$var wire 2 u& w [1:0] $end
$scope module M0 $end
$var wire 2 v& inputLines [1:0] $end
$var wire 1 w& outputLine $end
$var wire 1 x& selectLine $end
$var wire 1 y& w1 $end
$var wire 1 z& w2 $end
$var wire 1 {& w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 |& inputLines [1:0] $end
$var wire 1 }& outputLine $end
$var wire 1 ~& selectLine $end
$var wire 1 !' w1 $end
$var wire 1 "' w2 $end
$var wire 1 #' w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 $' inputLines [1:0] $end
$var wire 1 _& outputLine $end
$var wire 1 %' selectLine $end
$var wire 1 &' w1 $end
$var wire 1 '' w2 $end
$var wire 1 (' w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A12 $end
$var wire 1 )' Ainvert $end
$var wire 1 *' Binvert $end
$var wire 1 +' CarryIn $end
$var wire 1 ,' CarryOut $end
$var wire 1 -' Less $end
$var wire 2 .' Operation [1:0] $end
$var wire 1 /' Result $end
$var wire 1 0' a $end
$var wire 1 1' b $end
$var wire 2 2' mux0inputs [1:0] $end
$var wire 2 3' mux1inputs [1:0] $end
$var wire 4 4' mux2inputs [3:0] $end
$var wire 1 5' w1 $end
$var wire 1 6' w2 $end
$scope module P0 $end
$var wire 2 7' inputLines [1:0] $end
$var wire 1 5' outputLine $end
$var wire 1 )' selectLine $end
$var wire 1 8' w1 $end
$var wire 1 9' w2 $end
$var wire 1 :' w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 ;' inputLines [1:0] $end
$var wire 1 6' outputLine $end
$var wire 1 *' selectLine $end
$var wire 1 <' w1 $end
$var wire 1 =' w2 $end
$var wire 1 >' w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 5' a $end
$var wire 1 6' b $end
$var wire 1 +' cin $end
$var wire 1 ,' cout $end
$var wire 1 ?' sum $end
$var wire 1 @' w1 $end
$var wire 1 A' w2 $end
$var wire 1 B' w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 C' inputLines [3:0] $end
$var wire 1 /' outputLine $end
$var wire 2 D' selectLines [1:0] $end
$var wire 2 E' w [1:0] $end
$scope module M0 $end
$var wire 2 F' inputLines [1:0] $end
$var wire 1 G' outputLine $end
$var wire 1 H' selectLine $end
$var wire 1 I' w1 $end
$var wire 1 J' w2 $end
$var wire 1 K' w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 L' inputLines [1:0] $end
$var wire 1 M' outputLine $end
$var wire 1 N' selectLine $end
$var wire 1 O' w1 $end
$var wire 1 P' w2 $end
$var wire 1 Q' w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 R' inputLines [1:0] $end
$var wire 1 /' outputLine $end
$var wire 1 S' selectLine $end
$var wire 1 T' w1 $end
$var wire 1 U' w2 $end
$var wire 1 V' w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A13 $end
$var wire 1 W' Ainvert $end
$var wire 1 X' Binvert $end
$var wire 1 Y' CarryIn $end
$var wire 1 Z' CarryOut $end
$var wire 1 [' Less $end
$var wire 2 \' Operation [1:0] $end
$var wire 1 ]' Result $end
$var wire 1 ^' a $end
$var wire 1 _' b $end
$var wire 2 `' mux0inputs [1:0] $end
$var wire 2 a' mux1inputs [1:0] $end
$var wire 4 b' mux2inputs [3:0] $end
$var wire 1 c' w1 $end
$var wire 1 d' w2 $end
$scope module P0 $end
$var wire 2 e' inputLines [1:0] $end
$var wire 1 c' outputLine $end
$var wire 1 W' selectLine $end
$var wire 1 f' w1 $end
$var wire 1 g' w2 $end
$var wire 1 h' w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 i' inputLines [1:0] $end
$var wire 1 d' outputLine $end
$var wire 1 X' selectLine $end
$var wire 1 j' w1 $end
$var wire 1 k' w2 $end
$var wire 1 l' w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 c' a $end
$var wire 1 d' b $end
$var wire 1 Y' cin $end
$var wire 1 Z' cout $end
$var wire 1 m' sum $end
$var wire 1 n' w1 $end
$var wire 1 o' w2 $end
$var wire 1 p' w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 q' inputLines [3:0] $end
$var wire 1 ]' outputLine $end
$var wire 2 r' selectLines [1:0] $end
$var wire 2 s' w [1:0] $end
$scope module M0 $end
$var wire 2 t' inputLines [1:0] $end
$var wire 1 u' outputLine $end
$var wire 1 v' selectLine $end
$var wire 1 w' w1 $end
$var wire 1 x' w2 $end
$var wire 1 y' w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 z' inputLines [1:0] $end
$var wire 1 {' outputLine $end
$var wire 1 |' selectLine $end
$var wire 1 }' w1 $end
$var wire 1 ~' w2 $end
$var wire 1 !( w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 "( inputLines [1:0] $end
$var wire 1 ]' outputLine $end
$var wire 1 #( selectLine $end
$var wire 1 $( w1 $end
$var wire 1 %( w2 $end
$var wire 1 &( w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A14 $end
$var wire 1 '( Ainvert $end
$var wire 1 (( Binvert $end
$var wire 1 )( CarryIn $end
$var wire 1 *( CarryOut $end
$var wire 1 +( Less $end
$var wire 2 ,( Operation [1:0] $end
$var wire 1 -( Result $end
$var wire 1 .( a $end
$var wire 1 /( b $end
$var wire 2 0( mux0inputs [1:0] $end
$var wire 2 1( mux1inputs [1:0] $end
$var wire 4 2( mux2inputs [3:0] $end
$var wire 1 3( w1 $end
$var wire 1 4( w2 $end
$scope module P0 $end
$var wire 2 5( inputLines [1:0] $end
$var wire 1 3( outputLine $end
$var wire 1 '( selectLine $end
$var wire 1 6( w1 $end
$var wire 1 7( w2 $end
$var wire 1 8( w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 9( inputLines [1:0] $end
$var wire 1 4( outputLine $end
$var wire 1 (( selectLine $end
$var wire 1 :( w1 $end
$var wire 1 ;( w2 $end
$var wire 1 <( w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 3( a $end
$var wire 1 4( b $end
$var wire 1 )( cin $end
$var wire 1 *( cout $end
$var wire 1 =( sum $end
$var wire 1 >( w1 $end
$var wire 1 ?( w2 $end
$var wire 1 @( w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 A( inputLines [3:0] $end
$var wire 1 -( outputLine $end
$var wire 2 B( selectLines [1:0] $end
$var wire 2 C( w [1:0] $end
$scope module M0 $end
$var wire 2 D( inputLines [1:0] $end
$var wire 1 E( outputLine $end
$var wire 1 F( selectLine $end
$var wire 1 G( w1 $end
$var wire 1 H( w2 $end
$var wire 1 I( w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 J( inputLines [1:0] $end
$var wire 1 K( outputLine $end
$var wire 1 L( selectLine $end
$var wire 1 M( w1 $end
$var wire 1 N( w2 $end
$var wire 1 O( w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 P( inputLines [1:0] $end
$var wire 1 -( outputLine $end
$var wire 1 Q( selectLine $end
$var wire 1 R( w1 $end
$var wire 1 S( w2 $end
$var wire 1 T( w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A15 $end
$var wire 1 U( Ainvert $end
$var wire 1 V( Binvert $end
$var wire 1 W( CarryIn $end
$var wire 1 X( CarryOut $end
$var wire 1 Y( Less $end
$var wire 2 Z( Operation [1:0] $end
$var wire 1 [( Result $end
$var wire 1 \( a $end
$var wire 1 ]( b $end
$var wire 2 ^( mux0inputs [1:0] $end
$var wire 2 _( mux1inputs [1:0] $end
$var wire 4 `( mux2inputs [3:0] $end
$var wire 1 a( w1 $end
$var wire 1 b( w2 $end
$scope module P0 $end
$var wire 2 c( inputLines [1:0] $end
$var wire 1 a( outputLine $end
$var wire 1 U( selectLine $end
$var wire 1 d( w1 $end
$var wire 1 e( w2 $end
$var wire 1 f( w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 g( inputLines [1:0] $end
$var wire 1 b( outputLine $end
$var wire 1 V( selectLine $end
$var wire 1 h( w1 $end
$var wire 1 i( w2 $end
$var wire 1 j( w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 a( a $end
$var wire 1 b( b $end
$var wire 1 W( cin $end
$var wire 1 X( cout $end
$var wire 1 k( sum $end
$var wire 1 l( w1 $end
$var wire 1 m( w2 $end
$var wire 1 n( w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 o( inputLines [3:0] $end
$var wire 1 [( outputLine $end
$var wire 2 p( selectLines [1:0] $end
$var wire 2 q( w [1:0] $end
$scope module M0 $end
$var wire 2 r( inputLines [1:0] $end
$var wire 1 s( outputLine $end
$var wire 1 t( selectLine $end
$var wire 1 u( w1 $end
$var wire 1 v( w2 $end
$var wire 1 w( w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 x( inputLines [1:0] $end
$var wire 1 y( outputLine $end
$var wire 1 z( selectLine $end
$var wire 1 {( w1 $end
$var wire 1 |( w2 $end
$var wire 1 }( w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 ~( inputLines [1:0] $end
$var wire 1 [( outputLine $end
$var wire 1 !) selectLine $end
$var wire 1 ") w1 $end
$var wire 1 #) w2 $end
$var wire 1 $) w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A16 $end
$var wire 1 %) Ainvert $end
$var wire 1 &) Binvert $end
$var wire 1 ') CarryIn $end
$var wire 1 () CarryOut $end
$var wire 1 )) Less $end
$var wire 2 *) Operation [1:0] $end
$var wire 1 +) Result $end
$var wire 1 ,) a $end
$var wire 1 -) b $end
$var wire 2 .) mux0inputs [1:0] $end
$var wire 2 /) mux1inputs [1:0] $end
$var wire 4 0) mux2inputs [3:0] $end
$var wire 1 1) w1 $end
$var wire 1 2) w2 $end
$scope module P0 $end
$var wire 2 3) inputLines [1:0] $end
$var wire 1 1) outputLine $end
$var wire 1 %) selectLine $end
$var wire 1 4) w1 $end
$var wire 1 5) w2 $end
$var wire 1 6) w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 7) inputLines [1:0] $end
$var wire 1 2) outputLine $end
$var wire 1 &) selectLine $end
$var wire 1 8) w1 $end
$var wire 1 9) w2 $end
$var wire 1 :) w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 1) a $end
$var wire 1 2) b $end
$var wire 1 ') cin $end
$var wire 1 () cout $end
$var wire 1 ;) sum $end
$var wire 1 <) w1 $end
$var wire 1 =) w2 $end
$var wire 1 >) w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 ?) inputLines [3:0] $end
$var wire 1 +) outputLine $end
$var wire 2 @) selectLines [1:0] $end
$var wire 2 A) w [1:0] $end
$scope module M0 $end
$var wire 2 B) inputLines [1:0] $end
$var wire 1 C) outputLine $end
$var wire 1 D) selectLine $end
$var wire 1 E) w1 $end
$var wire 1 F) w2 $end
$var wire 1 G) w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 H) inputLines [1:0] $end
$var wire 1 I) outputLine $end
$var wire 1 J) selectLine $end
$var wire 1 K) w1 $end
$var wire 1 L) w2 $end
$var wire 1 M) w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 N) inputLines [1:0] $end
$var wire 1 +) outputLine $end
$var wire 1 O) selectLine $end
$var wire 1 P) w1 $end
$var wire 1 Q) w2 $end
$var wire 1 R) w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A17 $end
$var wire 1 S) Ainvert $end
$var wire 1 T) Binvert $end
$var wire 1 U) CarryIn $end
$var wire 1 V) CarryOut $end
$var wire 1 W) Less $end
$var wire 2 X) Operation [1:0] $end
$var wire 1 Y) Result $end
$var wire 1 Z) a $end
$var wire 1 [) b $end
$var wire 2 \) mux0inputs [1:0] $end
$var wire 2 ]) mux1inputs [1:0] $end
$var wire 4 ^) mux2inputs [3:0] $end
$var wire 1 _) w1 $end
$var wire 1 `) w2 $end
$scope module P0 $end
$var wire 2 a) inputLines [1:0] $end
$var wire 1 _) outputLine $end
$var wire 1 S) selectLine $end
$var wire 1 b) w1 $end
$var wire 1 c) w2 $end
$var wire 1 d) w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 e) inputLines [1:0] $end
$var wire 1 `) outputLine $end
$var wire 1 T) selectLine $end
$var wire 1 f) w1 $end
$var wire 1 g) w2 $end
$var wire 1 h) w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 _) a $end
$var wire 1 `) b $end
$var wire 1 U) cin $end
$var wire 1 V) cout $end
$var wire 1 i) sum $end
$var wire 1 j) w1 $end
$var wire 1 k) w2 $end
$var wire 1 l) w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 m) inputLines [3:0] $end
$var wire 1 Y) outputLine $end
$var wire 2 n) selectLines [1:0] $end
$var wire 2 o) w [1:0] $end
$scope module M0 $end
$var wire 2 p) inputLines [1:0] $end
$var wire 1 q) outputLine $end
$var wire 1 r) selectLine $end
$var wire 1 s) w1 $end
$var wire 1 t) w2 $end
$var wire 1 u) w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 v) inputLines [1:0] $end
$var wire 1 w) outputLine $end
$var wire 1 x) selectLine $end
$var wire 1 y) w1 $end
$var wire 1 z) w2 $end
$var wire 1 {) w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 |) inputLines [1:0] $end
$var wire 1 Y) outputLine $end
$var wire 1 }) selectLine $end
$var wire 1 ~) w1 $end
$var wire 1 !* w2 $end
$var wire 1 "* w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A18 $end
$var wire 1 #* Ainvert $end
$var wire 1 $* Binvert $end
$var wire 1 %* CarryIn $end
$var wire 1 &* CarryOut $end
$var wire 1 '* Less $end
$var wire 2 (* Operation [1:0] $end
$var wire 1 )* Result $end
$var wire 1 ** a $end
$var wire 1 +* b $end
$var wire 2 ,* mux0inputs [1:0] $end
$var wire 2 -* mux1inputs [1:0] $end
$var wire 4 .* mux2inputs [3:0] $end
$var wire 1 /* w1 $end
$var wire 1 0* w2 $end
$scope module P0 $end
$var wire 2 1* inputLines [1:0] $end
$var wire 1 /* outputLine $end
$var wire 1 #* selectLine $end
$var wire 1 2* w1 $end
$var wire 1 3* w2 $end
$var wire 1 4* w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 5* inputLines [1:0] $end
$var wire 1 0* outputLine $end
$var wire 1 $* selectLine $end
$var wire 1 6* w1 $end
$var wire 1 7* w2 $end
$var wire 1 8* w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 /* a $end
$var wire 1 0* b $end
$var wire 1 %* cin $end
$var wire 1 &* cout $end
$var wire 1 9* sum $end
$var wire 1 :* w1 $end
$var wire 1 ;* w2 $end
$var wire 1 <* w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 =* inputLines [3:0] $end
$var wire 1 )* outputLine $end
$var wire 2 >* selectLines [1:0] $end
$var wire 2 ?* w [1:0] $end
$scope module M0 $end
$var wire 2 @* inputLines [1:0] $end
$var wire 1 A* outputLine $end
$var wire 1 B* selectLine $end
$var wire 1 C* w1 $end
$var wire 1 D* w2 $end
$var wire 1 E* w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 F* inputLines [1:0] $end
$var wire 1 G* outputLine $end
$var wire 1 H* selectLine $end
$var wire 1 I* w1 $end
$var wire 1 J* w2 $end
$var wire 1 K* w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 L* inputLines [1:0] $end
$var wire 1 )* outputLine $end
$var wire 1 M* selectLine $end
$var wire 1 N* w1 $end
$var wire 1 O* w2 $end
$var wire 1 P* w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A19 $end
$var wire 1 Q* Ainvert $end
$var wire 1 R* Binvert $end
$var wire 1 S* CarryIn $end
$var wire 1 T* CarryOut $end
$var wire 1 U* Less $end
$var wire 2 V* Operation [1:0] $end
$var wire 1 W* Result $end
$var wire 1 X* a $end
$var wire 1 Y* b $end
$var wire 2 Z* mux0inputs [1:0] $end
$var wire 2 [* mux1inputs [1:0] $end
$var wire 4 \* mux2inputs [3:0] $end
$var wire 1 ]* w1 $end
$var wire 1 ^* w2 $end
$scope module P0 $end
$var wire 2 _* inputLines [1:0] $end
$var wire 1 ]* outputLine $end
$var wire 1 Q* selectLine $end
$var wire 1 `* w1 $end
$var wire 1 a* w2 $end
$var wire 1 b* w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 c* inputLines [1:0] $end
$var wire 1 ^* outputLine $end
$var wire 1 R* selectLine $end
$var wire 1 d* w1 $end
$var wire 1 e* w2 $end
$var wire 1 f* w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 ]* a $end
$var wire 1 ^* b $end
$var wire 1 S* cin $end
$var wire 1 T* cout $end
$var wire 1 g* sum $end
$var wire 1 h* w1 $end
$var wire 1 i* w2 $end
$var wire 1 j* w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 k* inputLines [3:0] $end
$var wire 1 W* outputLine $end
$var wire 2 l* selectLines [1:0] $end
$var wire 2 m* w [1:0] $end
$scope module M0 $end
$var wire 2 n* inputLines [1:0] $end
$var wire 1 o* outputLine $end
$var wire 1 p* selectLine $end
$var wire 1 q* w1 $end
$var wire 1 r* w2 $end
$var wire 1 s* w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 t* inputLines [1:0] $end
$var wire 1 u* outputLine $end
$var wire 1 v* selectLine $end
$var wire 1 w* w1 $end
$var wire 1 x* w2 $end
$var wire 1 y* w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 z* inputLines [1:0] $end
$var wire 1 W* outputLine $end
$var wire 1 {* selectLine $end
$var wire 1 |* w1 $end
$var wire 1 }* w2 $end
$var wire 1 ~* w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A20 $end
$var wire 1 !+ Ainvert $end
$var wire 1 "+ Binvert $end
$var wire 1 #+ CarryIn $end
$var wire 1 $+ CarryOut $end
$var wire 1 %+ Less $end
$var wire 2 &+ Operation [1:0] $end
$var wire 1 '+ Result $end
$var wire 1 (+ a $end
$var wire 1 )+ b $end
$var wire 2 *+ mux0inputs [1:0] $end
$var wire 2 ++ mux1inputs [1:0] $end
$var wire 4 ,+ mux2inputs [3:0] $end
$var wire 1 -+ w1 $end
$var wire 1 .+ w2 $end
$scope module P0 $end
$var wire 2 /+ inputLines [1:0] $end
$var wire 1 -+ outputLine $end
$var wire 1 !+ selectLine $end
$var wire 1 0+ w1 $end
$var wire 1 1+ w2 $end
$var wire 1 2+ w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 3+ inputLines [1:0] $end
$var wire 1 .+ outputLine $end
$var wire 1 "+ selectLine $end
$var wire 1 4+ w1 $end
$var wire 1 5+ w2 $end
$var wire 1 6+ w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 -+ a $end
$var wire 1 .+ b $end
$var wire 1 #+ cin $end
$var wire 1 $+ cout $end
$var wire 1 7+ sum $end
$var wire 1 8+ w1 $end
$var wire 1 9+ w2 $end
$var wire 1 :+ w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 ;+ inputLines [3:0] $end
$var wire 1 '+ outputLine $end
$var wire 2 <+ selectLines [1:0] $end
$var wire 2 =+ w [1:0] $end
$scope module M0 $end
$var wire 2 >+ inputLines [1:0] $end
$var wire 1 ?+ outputLine $end
$var wire 1 @+ selectLine $end
$var wire 1 A+ w1 $end
$var wire 1 B+ w2 $end
$var wire 1 C+ w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 D+ inputLines [1:0] $end
$var wire 1 E+ outputLine $end
$var wire 1 F+ selectLine $end
$var wire 1 G+ w1 $end
$var wire 1 H+ w2 $end
$var wire 1 I+ w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 J+ inputLines [1:0] $end
$var wire 1 '+ outputLine $end
$var wire 1 K+ selectLine $end
$var wire 1 L+ w1 $end
$var wire 1 M+ w2 $end
$var wire 1 N+ w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A21 $end
$var wire 1 O+ Ainvert $end
$var wire 1 P+ Binvert $end
$var wire 1 Q+ CarryIn $end
$var wire 1 R+ CarryOut $end
$var wire 1 S+ Less $end
$var wire 2 T+ Operation [1:0] $end
$var wire 1 U+ Result $end
$var wire 1 V+ a $end
$var wire 1 W+ b $end
$var wire 2 X+ mux0inputs [1:0] $end
$var wire 2 Y+ mux1inputs [1:0] $end
$var wire 4 Z+ mux2inputs [3:0] $end
$var wire 1 [+ w1 $end
$var wire 1 \+ w2 $end
$scope module P0 $end
$var wire 2 ]+ inputLines [1:0] $end
$var wire 1 [+ outputLine $end
$var wire 1 O+ selectLine $end
$var wire 1 ^+ w1 $end
$var wire 1 _+ w2 $end
$var wire 1 `+ w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 a+ inputLines [1:0] $end
$var wire 1 \+ outputLine $end
$var wire 1 P+ selectLine $end
$var wire 1 b+ w1 $end
$var wire 1 c+ w2 $end
$var wire 1 d+ w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 [+ a $end
$var wire 1 \+ b $end
$var wire 1 Q+ cin $end
$var wire 1 R+ cout $end
$var wire 1 e+ sum $end
$var wire 1 f+ w1 $end
$var wire 1 g+ w2 $end
$var wire 1 h+ w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 i+ inputLines [3:0] $end
$var wire 1 U+ outputLine $end
$var wire 2 j+ selectLines [1:0] $end
$var wire 2 k+ w [1:0] $end
$scope module M0 $end
$var wire 2 l+ inputLines [1:0] $end
$var wire 1 m+ outputLine $end
$var wire 1 n+ selectLine $end
$var wire 1 o+ w1 $end
$var wire 1 p+ w2 $end
$var wire 1 q+ w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 r+ inputLines [1:0] $end
$var wire 1 s+ outputLine $end
$var wire 1 t+ selectLine $end
$var wire 1 u+ w1 $end
$var wire 1 v+ w2 $end
$var wire 1 w+ w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 x+ inputLines [1:0] $end
$var wire 1 U+ outputLine $end
$var wire 1 y+ selectLine $end
$var wire 1 z+ w1 $end
$var wire 1 {+ w2 $end
$var wire 1 |+ w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A22 $end
$var wire 1 }+ Ainvert $end
$var wire 1 ~+ Binvert $end
$var wire 1 !, CarryIn $end
$var wire 1 ", CarryOut $end
$var wire 1 #, Less $end
$var wire 2 $, Operation [1:0] $end
$var wire 1 %, Result $end
$var wire 1 &, a $end
$var wire 1 ', b $end
$var wire 2 (, mux0inputs [1:0] $end
$var wire 2 ), mux1inputs [1:0] $end
$var wire 4 *, mux2inputs [3:0] $end
$var wire 1 +, w1 $end
$var wire 1 ,, w2 $end
$scope module P0 $end
$var wire 2 -, inputLines [1:0] $end
$var wire 1 +, outputLine $end
$var wire 1 }+ selectLine $end
$var wire 1 ., w1 $end
$var wire 1 /, w2 $end
$var wire 1 0, w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 1, inputLines [1:0] $end
$var wire 1 ,, outputLine $end
$var wire 1 ~+ selectLine $end
$var wire 1 2, w1 $end
$var wire 1 3, w2 $end
$var wire 1 4, w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 +, a $end
$var wire 1 ,, b $end
$var wire 1 !, cin $end
$var wire 1 ", cout $end
$var wire 1 5, sum $end
$var wire 1 6, w1 $end
$var wire 1 7, w2 $end
$var wire 1 8, w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 9, inputLines [3:0] $end
$var wire 1 %, outputLine $end
$var wire 2 :, selectLines [1:0] $end
$var wire 2 ;, w [1:0] $end
$scope module M0 $end
$var wire 2 <, inputLines [1:0] $end
$var wire 1 =, outputLine $end
$var wire 1 >, selectLine $end
$var wire 1 ?, w1 $end
$var wire 1 @, w2 $end
$var wire 1 A, w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 B, inputLines [1:0] $end
$var wire 1 C, outputLine $end
$var wire 1 D, selectLine $end
$var wire 1 E, w1 $end
$var wire 1 F, w2 $end
$var wire 1 G, w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 H, inputLines [1:0] $end
$var wire 1 %, outputLine $end
$var wire 1 I, selectLine $end
$var wire 1 J, w1 $end
$var wire 1 K, w2 $end
$var wire 1 L, w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A23 $end
$var wire 1 M, Ainvert $end
$var wire 1 N, Binvert $end
$var wire 1 O, CarryIn $end
$var wire 1 P, CarryOut $end
$var wire 1 Q, Less $end
$var wire 2 R, Operation [1:0] $end
$var wire 1 S, Result $end
$var wire 1 T, a $end
$var wire 1 U, b $end
$var wire 2 V, mux0inputs [1:0] $end
$var wire 2 W, mux1inputs [1:0] $end
$var wire 4 X, mux2inputs [3:0] $end
$var wire 1 Y, w1 $end
$var wire 1 Z, w2 $end
$scope module P0 $end
$var wire 2 [, inputLines [1:0] $end
$var wire 1 Y, outputLine $end
$var wire 1 M, selectLine $end
$var wire 1 \, w1 $end
$var wire 1 ], w2 $end
$var wire 1 ^, w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 _, inputLines [1:0] $end
$var wire 1 Z, outputLine $end
$var wire 1 N, selectLine $end
$var wire 1 `, w1 $end
$var wire 1 a, w2 $end
$var wire 1 b, w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 Y, a $end
$var wire 1 Z, b $end
$var wire 1 O, cin $end
$var wire 1 P, cout $end
$var wire 1 c, sum $end
$var wire 1 d, w1 $end
$var wire 1 e, w2 $end
$var wire 1 f, w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 g, inputLines [3:0] $end
$var wire 1 S, outputLine $end
$var wire 2 h, selectLines [1:0] $end
$var wire 2 i, w [1:0] $end
$scope module M0 $end
$var wire 2 j, inputLines [1:0] $end
$var wire 1 k, outputLine $end
$var wire 1 l, selectLine $end
$var wire 1 m, w1 $end
$var wire 1 n, w2 $end
$var wire 1 o, w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 p, inputLines [1:0] $end
$var wire 1 q, outputLine $end
$var wire 1 r, selectLine $end
$var wire 1 s, w1 $end
$var wire 1 t, w2 $end
$var wire 1 u, w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 v, inputLines [1:0] $end
$var wire 1 S, outputLine $end
$var wire 1 w, selectLine $end
$var wire 1 x, w1 $end
$var wire 1 y, w2 $end
$var wire 1 z, w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A24 $end
$var wire 1 {, Ainvert $end
$var wire 1 |, Binvert $end
$var wire 1 }, CarryIn $end
$var wire 1 ~, CarryOut $end
$var wire 1 !- Less $end
$var wire 2 "- Operation [1:0] $end
$var wire 1 #- Result $end
$var wire 1 $- a $end
$var wire 1 %- b $end
$var wire 2 &- mux0inputs [1:0] $end
$var wire 2 '- mux1inputs [1:0] $end
$var wire 4 (- mux2inputs [3:0] $end
$var wire 1 )- w1 $end
$var wire 1 *- w2 $end
$scope module P0 $end
$var wire 2 +- inputLines [1:0] $end
$var wire 1 )- outputLine $end
$var wire 1 {, selectLine $end
$var wire 1 ,- w1 $end
$var wire 1 -- w2 $end
$var wire 1 .- w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 /- inputLines [1:0] $end
$var wire 1 *- outputLine $end
$var wire 1 |, selectLine $end
$var wire 1 0- w1 $end
$var wire 1 1- w2 $end
$var wire 1 2- w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 )- a $end
$var wire 1 *- b $end
$var wire 1 }, cin $end
$var wire 1 ~, cout $end
$var wire 1 3- sum $end
$var wire 1 4- w1 $end
$var wire 1 5- w2 $end
$var wire 1 6- w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 7- inputLines [3:0] $end
$var wire 1 #- outputLine $end
$var wire 2 8- selectLines [1:0] $end
$var wire 2 9- w [1:0] $end
$scope module M0 $end
$var wire 2 :- inputLines [1:0] $end
$var wire 1 ;- outputLine $end
$var wire 1 <- selectLine $end
$var wire 1 =- w1 $end
$var wire 1 >- w2 $end
$var wire 1 ?- w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 @- inputLines [1:0] $end
$var wire 1 A- outputLine $end
$var wire 1 B- selectLine $end
$var wire 1 C- w1 $end
$var wire 1 D- w2 $end
$var wire 1 E- w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 F- inputLines [1:0] $end
$var wire 1 #- outputLine $end
$var wire 1 G- selectLine $end
$var wire 1 H- w1 $end
$var wire 1 I- w2 $end
$var wire 1 J- w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A25 $end
$var wire 1 K- Ainvert $end
$var wire 1 L- Binvert $end
$var wire 1 M- CarryIn $end
$var wire 1 N- CarryOut $end
$var wire 1 O- Less $end
$var wire 2 P- Operation [1:0] $end
$var wire 1 Q- Result $end
$var wire 1 R- a $end
$var wire 1 S- b $end
$var wire 2 T- mux0inputs [1:0] $end
$var wire 2 U- mux1inputs [1:0] $end
$var wire 4 V- mux2inputs [3:0] $end
$var wire 1 W- w1 $end
$var wire 1 X- w2 $end
$scope module P0 $end
$var wire 2 Y- inputLines [1:0] $end
$var wire 1 W- outputLine $end
$var wire 1 K- selectLine $end
$var wire 1 Z- w1 $end
$var wire 1 [- w2 $end
$var wire 1 \- w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 ]- inputLines [1:0] $end
$var wire 1 X- outputLine $end
$var wire 1 L- selectLine $end
$var wire 1 ^- w1 $end
$var wire 1 _- w2 $end
$var wire 1 `- w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 W- a $end
$var wire 1 X- b $end
$var wire 1 M- cin $end
$var wire 1 N- cout $end
$var wire 1 a- sum $end
$var wire 1 b- w1 $end
$var wire 1 c- w2 $end
$var wire 1 d- w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 e- inputLines [3:0] $end
$var wire 1 Q- outputLine $end
$var wire 2 f- selectLines [1:0] $end
$var wire 2 g- w [1:0] $end
$scope module M0 $end
$var wire 2 h- inputLines [1:0] $end
$var wire 1 i- outputLine $end
$var wire 1 j- selectLine $end
$var wire 1 k- w1 $end
$var wire 1 l- w2 $end
$var wire 1 m- w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 n- inputLines [1:0] $end
$var wire 1 o- outputLine $end
$var wire 1 p- selectLine $end
$var wire 1 q- w1 $end
$var wire 1 r- w2 $end
$var wire 1 s- w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 t- inputLines [1:0] $end
$var wire 1 Q- outputLine $end
$var wire 1 u- selectLine $end
$var wire 1 v- w1 $end
$var wire 1 w- w2 $end
$var wire 1 x- w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A26 $end
$var wire 1 y- Ainvert $end
$var wire 1 z- Binvert $end
$var wire 1 {- CarryIn $end
$var wire 1 |- CarryOut $end
$var wire 1 }- Less $end
$var wire 2 ~- Operation [1:0] $end
$var wire 1 !. Result $end
$var wire 1 ". a $end
$var wire 1 #. b $end
$var wire 2 $. mux0inputs [1:0] $end
$var wire 2 %. mux1inputs [1:0] $end
$var wire 4 &. mux2inputs [3:0] $end
$var wire 1 '. w1 $end
$var wire 1 (. w2 $end
$scope module P0 $end
$var wire 2 ). inputLines [1:0] $end
$var wire 1 '. outputLine $end
$var wire 1 y- selectLine $end
$var wire 1 *. w1 $end
$var wire 1 +. w2 $end
$var wire 1 ,. w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 -. inputLines [1:0] $end
$var wire 1 (. outputLine $end
$var wire 1 z- selectLine $end
$var wire 1 .. w1 $end
$var wire 1 /. w2 $end
$var wire 1 0. w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 '. a $end
$var wire 1 (. b $end
$var wire 1 {- cin $end
$var wire 1 |- cout $end
$var wire 1 1. sum $end
$var wire 1 2. w1 $end
$var wire 1 3. w2 $end
$var wire 1 4. w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 5. inputLines [3:0] $end
$var wire 1 !. outputLine $end
$var wire 2 6. selectLines [1:0] $end
$var wire 2 7. w [1:0] $end
$scope module M0 $end
$var wire 2 8. inputLines [1:0] $end
$var wire 1 9. outputLine $end
$var wire 1 :. selectLine $end
$var wire 1 ;. w1 $end
$var wire 1 <. w2 $end
$var wire 1 =. w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 >. inputLines [1:0] $end
$var wire 1 ?. outputLine $end
$var wire 1 @. selectLine $end
$var wire 1 A. w1 $end
$var wire 1 B. w2 $end
$var wire 1 C. w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 D. inputLines [1:0] $end
$var wire 1 !. outputLine $end
$var wire 1 E. selectLine $end
$var wire 1 F. w1 $end
$var wire 1 G. w2 $end
$var wire 1 H. w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A27 $end
$var wire 1 I. Ainvert $end
$var wire 1 J. Binvert $end
$var wire 1 K. CarryIn $end
$var wire 1 L. CarryOut $end
$var wire 1 M. Less $end
$var wire 2 N. Operation [1:0] $end
$var wire 1 O. Result $end
$var wire 1 P. a $end
$var wire 1 Q. b $end
$var wire 2 R. mux0inputs [1:0] $end
$var wire 2 S. mux1inputs [1:0] $end
$var wire 4 T. mux2inputs [3:0] $end
$var wire 1 U. w1 $end
$var wire 1 V. w2 $end
$scope module P0 $end
$var wire 2 W. inputLines [1:0] $end
$var wire 1 U. outputLine $end
$var wire 1 I. selectLine $end
$var wire 1 X. w1 $end
$var wire 1 Y. w2 $end
$var wire 1 Z. w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 [. inputLines [1:0] $end
$var wire 1 V. outputLine $end
$var wire 1 J. selectLine $end
$var wire 1 \. w1 $end
$var wire 1 ]. w2 $end
$var wire 1 ^. w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 U. a $end
$var wire 1 V. b $end
$var wire 1 K. cin $end
$var wire 1 L. cout $end
$var wire 1 _. sum $end
$var wire 1 `. w1 $end
$var wire 1 a. w2 $end
$var wire 1 b. w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 c. inputLines [3:0] $end
$var wire 1 O. outputLine $end
$var wire 2 d. selectLines [1:0] $end
$var wire 2 e. w [1:0] $end
$scope module M0 $end
$var wire 2 f. inputLines [1:0] $end
$var wire 1 g. outputLine $end
$var wire 1 h. selectLine $end
$var wire 1 i. w1 $end
$var wire 1 j. w2 $end
$var wire 1 k. w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 l. inputLines [1:0] $end
$var wire 1 m. outputLine $end
$var wire 1 n. selectLine $end
$var wire 1 o. w1 $end
$var wire 1 p. w2 $end
$var wire 1 q. w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 r. inputLines [1:0] $end
$var wire 1 O. outputLine $end
$var wire 1 s. selectLine $end
$var wire 1 t. w1 $end
$var wire 1 u. w2 $end
$var wire 1 v. w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A28 $end
$var wire 1 w. Ainvert $end
$var wire 1 x. Binvert $end
$var wire 1 y. CarryIn $end
$var wire 1 z. CarryOut $end
$var wire 1 {. Less $end
$var wire 2 |. Operation [1:0] $end
$var wire 1 }. Result $end
$var wire 1 ~. a $end
$var wire 1 !/ b $end
$var wire 2 "/ mux0inputs [1:0] $end
$var wire 2 #/ mux1inputs [1:0] $end
$var wire 4 $/ mux2inputs [3:0] $end
$var wire 1 %/ w1 $end
$var wire 1 &/ w2 $end
$scope module P0 $end
$var wire 2 '/ inputLines [1:0] $end
$var wire 1 %/ outputLine $end
$var wire 1 w. selectLine $end
$var wire 1 (/ w1 $end
$var wire 1 )/ w2 $end
$var wire 1 */ w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 +/ inputLines [1:0] $end
$var wire 1 &/ outputLine $end
$var wire 1 x. selectLine $end
$var wire 1 ,/ w1 $end
$var wire 1 -/ w2 $end
$var wire 1 ./ w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 %/ a $end
$var wire 1 &/ b $end
$var wire 1 y. cin $end
$var wire 1 z. cout $end
$var wire 1 // sum $end
$var wire 1 0/ w1 $end
$var wire 1 1/ w2 $end
$var wire 1 2/ w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 3/ inputLines [3:0] $end
$var wire 1 }. outputLine $end
$var wire 2 4/ selectLines [1:0] $end
$var wire 2 5/ w [1:0] $end
$scope module M0 $end
$var wire 2 6/ inputLines [1:0] $end
$var wire 1 7/ outputLine $end
$var wire 1 8/ selectLine $end
$var wire 1 9/ w1 $end
$var wire 1 :/ w2 $end
$var wire 1 ;/ w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 </ inputLines [1:0] $end
$var wire 1 =/ outputLine $end
$var wire 1 >/ selectLine $end
$var wire 1 ?/ w1 $end
$var wire 1 @/ w2 $end
$var wire 1 A/ w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 B/ inputLines [1:0] $end
$var wire 1 }. outputLine $end
$var wire 1 C/ selectLine $end
$var wire 1 D/ w1 $end
$var wire 1 E/ w2 $end
$var wire 1 F/ w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A29 $end
$var wire 1 G/ Ainvert $end
$var wire 1 H/ Binvert $end
$var wire 1 I/ CarryIn $end
$var wire 1 J/ CarryOut $end
$var wire 1 K/ Less $end
$var wire 2 L/ Operation [1:0] $end
$var wire 1 M/ Result $end
$var wire 1 N/ a $end
$var wire 1 O/ b $end
$var wire 2 P/ mux0inputs [1:0] $end
$var wire 2 Q/ mux1inputs [1:0] $end
$var wire 4 R/ mux2inputs [3:0] $end
$var wire 1 S/ w1 $end
$var wire 1 T/ w2 $end
$scope module P0 $end
$var wire 2 U/ inputLines [1:0] $end
$var wire 1 S/ outputLine $end
$var wire 1 G/ selectLine $end
$var wire 1 V/ w1 $end
$var wire 1 W/ w2 $end
$var wire 1 X/ w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 Y/ inputLines [1:0] $end
$var wire 1 T/ outputLine $end
$var wire 1 H/ selectLine $end
$var wire 1 Z/ w1 $end
$var wire 1 [/ w2 $end
$var wire 1 \/ w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 S/ a $end
$var wire 1 T/ b $end
$var wire 1 I/ cin $end
$var wire 1 J/ cout $end
$var wire 1 ]/ sum $end
$var wire 1 ^/ w1 $end
$var wire 1 _/ w2 $end
$var wire 1 `/ w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 a/ inputLines [3:0] $end
$var wire 1 M/ outputLine $end
$var wire 2 b/ selectLines [1:0] $end
$var wire 2 c/ w [1:0] $end
$scope module M0 $end
$var wire 2 d/ inputLines [1:0] $end
$var wire 1 e/ outputLine $end
$var wire 1 f/ selectLine $end
$var wire 1 g/ w1 $end
$var wire 1 h/ w2 $end
$var wire 1 i/ w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 j/ inputLines [1:0] $end
$var wire 1 k/ outputLine $end
$var wire 1 l/ selectLine $end
$var wire 1 m/ w1 $end
$var wire 1 n/ w2 $end
$var wire 1 o/ w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 p/ inputLines [1:0] $end
$var wire 1 M/ outputLine $end
$var wire 1 q/ selectLine $end
$var wire 1 r/ w1 $end
$var wire 1 s/ w2 $end
$var wire 1 t/ w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A30 $end
$var wire 1 u/ Ainvert $end
$var wire 1 v/ Binvert $end
$var wire 1 w/ CarryIn $end
$var wire 1 x/ CarryOut $end
$var wire 1 y/ Less $end
$var wire 2 z/ Operation [1:0] $end
$var wire 1 {/ Result $end
$var wire 1 |/ a $end
$var wire 1 }/ b $end
$var wire 2 ~/ mux0inputs [1:0] $end
$var wire 2 !0 mux1inputs [1:0] $end
$var wire 4 "0 mux2inputs [3:0] $end
$var wire 1 #0 w1 $end
$var wire 1 $0 w2 $end
$scope module P0 $end
$var wire 2 %0 inputLines [1:0] $end
$var wire 1 #0 outputLine $end
$var wire 1 u/ selectLine $end
$var wire 1 &0 w1 $end
$var wire 1 '0 w2 $end
$var wire 1 (0 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 )0 inputLines [1:0] $end
$var wire 1 $0 outputLine $end
$var wire 1 v/ selectLine $end
$var wire 1 *0 w1 $end
$var wire 1 +0 w2 $end
$var wire 1 ,0 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 #0 a $end
$var wire 1 $0 b $end
$var wire 1 w/ cin $end
$var wire 1 x/ cout $end
$var wire 1 -0 sum $end
$var wire 1 .0 w1 $end
$var wire 1 /0 w2 $end
$var wire 1 00 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 10 inputLines [3:0] $end
$var wire 1 {/ outputLine $end
$var wire 2 20 selectLines [1:0] $end
$var wire 2 30 w [1:0] $end
$scope module M0 $end
$var wire 2 40 inputLines [1:0] $end
$var wire 1 50 outputLine $end
$var wire 1 60 selectLine $end
$var wire 1 70 w1 $end
$var wire 1 80 w2 $end
$var wire 1 90 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 :0 inputLines [1:0] $end
$var wire 1 ;0 outputLine $end
$var wire 1 <0 selectLine $end
$var wire 1 =0 w1 $end
$var wire 1 >0 w2 $end
$var wire 1 ?0 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 @0 inputLines [1:0] $end
$var wire 1 {/ outputLine $end
$var wire 1 A0 selectLine $end
$var wire 1 B0 w1 $end
$var wire 1 C0 w2 $end
$var wire 1 D0 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A31 $end
$var wire 1 E0 Ainvert $end
$var wire 1 F0 Binvert $end
$var wire 1 G0 CarryIn $end
$var wire 1 H0 CarryOut $end
$var wire 1 I0 Less $end
$var wire 2 J0 Operation [1:0] $end
$var wire 1 K0 Result $end
$var wire 1 L0 a $end
$var wire 1 M0 b $end
$var wire 2 N0 mux0inputs [1:0] $end
$var wire 2 O0 mux1inputs [1:0] $end
$var wire 4 P0 mux2inputs [3:0] $end
$var wire 1 Q0 w1 $end
$var wire 1 R0 w2 $end
$scope module P0 $end
$var wire 2 S0 inputLines [1:0] $end
$var wire 1 Q0 outputLine $end
$var wire 1 E0 selectLine $end
$var wire 1 T0 w1 $end
$var wire 1 U0 w2 $end
$var wire 1 V0 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 W0 inputLines [1:0] $end
$var wire 1 R0 outputLine $end
$var wire 1 F0 selectLine $end
$var wire 1 X0 w1 $end
$var wire 1 Y0 w2 $end
$var wire 1 Z0 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 Q0 a $end
$var wire 1 R0 b $end
$var wire 1 G0 cin $end
$var wire 1 H0 cout $end
$var wire 1 [0 sum $end
$var wire 1 \0 w1 $end
$var wire 1 ]0 w2 $end
$var wire 1 ^0 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 _0 inputLines [3:0] $end
$var wire 1 K0 outputLine $end
$var wire 2 `0 selectLines [1:0] $end
$var wire 2 a0 w [1:0] $end
$scope module M0 $end
$var wire 2 b0 inputLines [1:0] $end
$var wire 1 c0 outputLine $end
$var wire 1 d0 selectLine $end
$var wire 1 e0 w1 $end
$var wire 1 f0 w2 $end
$var wire 1 g0 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 h0 inputLines [1:0] $end
$var wire 1 i0 outputLine $end
$var wire 1 j0 selectLine $end
$var wire 1 k0 w1 $end
$var wire 1 l0 w2 $end
$var wire 1 m0 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 n0 inputLines [1:0] $end
$var wire 1 K0 outputLine $end
$var wire 1 o0 selectLine $end
$var wire 1 p0 w1 $end
$var wire 1 q0 w2 $end
$var wire 1 r0 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A32 $end
$var wire 1 s0 Ainvert $end
$var wire 1 t0 Binvert $end
$var wire 1 u0 CarryIn $end
$var wire 1 v0 CarryOut $end
$var wire 1 w0 Less $end
$var wire 2 x0 Operation [1:0] $end
$var wire 1 y0 Result $end
$var wire 1 z0 a $end
$var wire 1 {0 b $end
$var wire 2 |0 mux0inputs [1:0] $end
$var wire 2 }0 mux1inputs [1:0] $end
$var wire 4 ~0 mux2inputs [3:0] $end
$var wire 1 !1 w1 $end
$var wire 1 "1 w2 $end
$scope module P0 $end
$var wire 2 #1 inputLines [1:0] $end
$var wire 1 !1 outputLine $end
$var wire 1 s0 selectLine $end
$var wire 1 $1 w1 $end
$var wire 1 %1 w2 $end
$var wire 1 &1 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 '1 inputLines [1:0] $end
$var wire 1 "1 outputLine $end
$var wire 1 t0 selectLine $end
$var wire 1 (1 w1 $end
$var wire 1 )1 w2 $end
$var wire 1 *1 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 !1 a $end
$var wire 1 "1 b $end
$var wire 1 u0 cin $end
$var wire 1 v0 cout $end
$var wire 1 +1 sum $end
$var wire 1 ,1 w1 $end
$var wire 1 -1 w2 $end
$var wire 1 .1 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 /1 inputLines [3:0] $end
$var wire 1 y0 outputLine $end
$var wire 2 01 selectLines [1:0] $end
$var wire 2 11 w [1:0] $end
$scope module M0 $end
$var wire 2 21 inputLines [1:0] $end
$var wire 1 31 outputLine $end
$var wire 1 41 selectLine $end
$var wire 1 51 w1 $end
$var wire 1 61 w2 $end
$var wire 1 71 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 81 inputLines [1:0] $end
$var wire 1 91 outputLine $end
$var wire 1 :1 selectLine $end
$var wire 1 ;1 w1 $end
$var wire 1 <1 w2 $end
$var wire 1 =1 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 >1 inputLines [1:0] $end
$var wire 1 y0 outputLine $end
$var wire 1 ?1 selectLine $end
$var wire 1 @1 w1 $end
$var wire 1 A1 w2 $end
$var wire 1 B1 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A33 $end
$var wire 1 C1 Ainvert $end
$var wire 1 D1 Binvert $end
$var wire 1 E1 CarryIn $end
$var wire 1 F1 CarryOut $end
$var wire 1 G1 Less $end
$var wire 2 H1 Operation [1:0] $end
$var wire 1 I1 Result $end
$var wire 1 J1 a $end
$var wire 1 K1 b $end
$var wire 2 L1 mux0inputs [1:0] $end
$var wire 2 M1 mux1inputs [1:0] $end
$var wire 4 N1 mux2inputs [3:0] $end
$var wire 1 O1 w1 $end
$var wire 1 P1 w2 $end
$scope module P0 $end
$var wire 2 Q1 inputLines [1:0] $end
$var wire 1 O1 outputLine $end
$var wire 1 C1 selectLine $end
$var wire 1 R1 w1 $end
$var wire 1 S1 w2 $end
$var wire 1 T1 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 U1 inputLines [1:0] $end
$var wire 1 P1 outputLine $end
$var wire 1 D1 selectLine $end
$var wire 1 V1 w1 $end
$var wire 1 W1 w2 $end
$var wire 1 X1 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 O1 a $end
$var wire 1 P1 b $end
$var wire 1 E1 cin $end
$var wire 1 F1 cout $end
$var wire 1 Y1 sum $end
$var wire 1 Z1 w1 $end
$var wire 1 [1 w2 $end
$var wire 1 \1 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 ]1 inputLines [3:0] $end
$var wire 1 I1 outputLine $end
$var wire 2 ^1 selectLines [1:0] $end
$var wire 2 _1 w [1:0] $end
$scope module M0 $end
$var wire 2 `1 inputLines [1:0] $end
$var wire 1 a1 outputLine $end
$var wire 1 b1 selectLine $end
$var wire 1 c1 w1 $end
$var wire 1 d1 w2 $end
$var wire 1 e1 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 f1 inputLines [1:0] $end
$var wire 1 g1 outputLine $end
$var wire 1 h1 selectLine $end
$var wire 1 i1 w1 $end
$var wire 1 j1 w2 $end
$var wire 1 k1 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 l1 inputLines [1:0] $end
$var wire 1 I1 outputLine $end
$var wire 1 m1 selectLine $end
$var wire 1 n1 w1 $end
$var wire 1 o1 w2 $end
$var wire 1 p1 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A34 $end
$var wire 1 q1 Ainvert $end
$var wire 1 r1 Binvert $end
$var wire 1 s1 CarryIn $end
$var wire 1 t1 CarryOut $end
$var wire 1 u1 Less $end
$var wire 2 v1 Operation [1:0] $end
$var wire 1 w1 Result $end
$var wire 1 x1 a $end
$var wire 1 y1 b $end
$var wire 2 z1 mux0inputs [1:0] $end
$var wire 2 {1 mux1inputs [1:0] $end
$var wire 4 |1 mux2inputs [3:0] $end
$var wire 1 }1 w1 $end
$var wire 1 ~1 w2 $end
$scope module P0 $end
$var wire 2 !2 inputLines [1:0] $end
$var wire 1 }1 outputLine $end
$var wire 1 q1 selectLine $end
$var wire 1 "2 w1 $end
$var wire 1 #2 w2 $end
$var wire 1 $2 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 %2 inputLines [1:0] $end
$var wire 1 ~1 outputLine $end
$var wire 1 r1 selectLine $end
$var wire 1 &2 w1 $end
$var wire 1 '2 w2 $end
$var wire 1 (2 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 }1 a $end
$var wire 1 ~1 b $end
$var wire 1 s1 cin $end
$var wire 1 t1 cout $end
$var wire 1 )2 sum $end
$var wire 1 *2 w1 $end
$var wire 1 +2 w2 $end
$var wire 1 ,2 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 -2 inputLines [3:0] $end
$var wire 1 w1 outputLine $end
$var wire 2 .2 selectLines [1:0] $end
$var wire 2 /2 w [1:0] $end
$scope module M0 $end
$var wire 2 02 inputLines [1:0] $end
$var wire 1 12 outputLine $end
$var wire 1 22 selectLine $end
$var wire 1 32 w1 $end
$var wire 1 42 w2 $end
$var wire 1 52 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 62 inputLines [1:0] $end
$var wire 1 72 outputLine $end
$var wire 1 82 selectLine $end
$var wire 1 92 w1 $end
$var wire 1 :2 w2 $end
$var wire 1 ;2 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 <2 inputLines [1:0] $end
$var wire 1 w1 outputLine $end
$var wire 1 =2 selectLine $end
$var wire 1 >2 w1 $end
$var wire 1 ?2 w2 $end
$var wire 1 @2 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A35 $end
$var wire 1 A2 Ainvert $end
$var wire 1 B2 Binvert $end
$var wire 1 C2 CarryIn $end
$var wire 1 D2 CarryOut $end
$var wire 1 E2 Less $end
$var wire 2 F2 Operation [1:0] $end
$var wire 1 G2 Result $end
$var wire 1 H2 a $end
$var wire 1 I2 b $end
$var wire 2 J2 mux0inputs [1:0] $end
$var wire 2 K2 mux1inputs [1:0] $end
$var wire 4 L2 mux2inputs [3:0] $end
$var wire 1 M2 w1 $end
$var wire 1 N2 w2 $end
$scope module P0 $end
$var wire 2 O2 inputLines [1:0] $end
$var wire 1 M2 outputLine $end
$var wire 1 A2 selectLine $end
$var wire 1 P2 w1 $end
$var wire 1 Q2 w2 $end
$var wire 1 R2 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 S2 inputLines [1:0] $end
$var wire 1 N2 outputLine $end
$var wire 1 B2 selectLine $end
$var wire 1 T2 w1 $end
$var wire 1 U2 w2 $end
$var wire 1 V2 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 M2 a $end
$var wire 1 N2 b $end
$var wire 1 C2 cin $end
$var wire 1 D2 cout $end
$var wire 1 W2 sum $end
$var wire 1 X2 w1 $end
$var wire 1 Y2 w2 $end
$var wire 1 Z2 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 [2 inputLines [3:0] $end
$var wire 1 G2 outputLine $end
$var wire 2 \2 selectLines [1:0] $end
$var wire 2 ]2 w [1:0] $end
$scope module M0 $end
$var wire 2 ^2 inputLines [1:0] $end
$var wire 1 _2 outputLine $end
$var wire 1 `2 selectLine $end
$var wire 1 a2 w1 $end
$var wire 1 b2 w2 $end
$var wire 1 c2 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 d2 inputLines [1:0] $end
$var wire 1 e2 outputLine $end
$var wire 1 f2 selectLine $end
$var wire 1 g2 w1 $end
$var wire 1 h2 w2 $end
$var wire 1 i2 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 j2 inputLines [1:0] $end
$var wire 1 G2 outputLine $end
$var wire 1 k2 selectLine $end
$var wire 1 l2 w1 $end
$var wire 1 m2 w2 $end
$var wire 1 n2 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A36 $end
$var wire 1 o2 Ainvert $end
$var wire 1 p2 Binvert $end
$var wire 1 q2 CarryIn $end
$var wire 1 r2 CarryOut $end
$var wire 1 s2 Less $end
$var wire 2 t2 Operation [1:0] $end
$var wire 1 u2 Result $end
$var wire 1 v2 a $end
$var wire 1 w2 b $end
$var wire 2 x2 mux0inputs [1:0] $end
$var wire 2 y2 mux1inputs [1:0] $end
$var wire 4 z2 mux2inputs [3:0] $end
$var wire 1 {2 w1 $end
$var wire 1 |2 w2 $end
$scope module P0 $end
$var wire 2 }2 inputLines [1:0] $end
$var wire 1 {2 outputLine $end
$var wire 1 o2 selectLine $end
$var wire 1 ~2 w1 $end
$var wire 1 !3 w2 $end
$var wire 1 "3 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 #3 inputLines [1:0] $end
$var wire 1 |2 outputLine $end
$var wire 1 p2 selectLine $end
$var wire 1 $3 w1 $end
$var wire 1 %3 w2 $end
$var wire 1 &3 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 {2 a $end
$var wire 1 |2 b $end
$var wire 1 q2 cin $end
$var wire 1 r2 cout $end
$var wire 1 '3 sum $end
$var wire 1 (3 w1 $end
$var wire 1 )3 w2 $end
$var wire 1 *3 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 +3 inputLines [3:0] $end
$var wire 1 u2 outputLine $end
$var wire 2 ,3 selectLines [1:0] $end
$var wire 2 -3 w [1:0] $end
$scope module M0 $end
$var wire 2 .3 inputLines [1:0] $end
$var wire 1 /3 outputLine $end
$var wire 1 03 selectLine $end
$var wire 1 13 w1 $end
$var wire 1 23 w2 $end
$var wire 1 33 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 43 inputLines [1:0] $end
$var wire 1 53 outputLine $end
$var wire 1 63 selectLine $end
$var wire 1 73 w1 $end
$var wire 1 83 w2 $end
$var wire 1 93 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 :3 inputLines [1:0] $end
$var wire 1 u2 outputLine $end
$var wire 1 ;3 selectLine $end
$var wire 1 <3 w1 $end
$var wire 1 =3 w2 $end
$var wire 1 >3 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A37 $end
$var wire 1 ?3 Ainvert $end
$var wire 1 @3 Binvert $end
$var wire 1 A3 CarryIn $end
$var wire 1 B3 CarryOut $end
$var wire 1 C3 Less $end
$var wire 2 D3 Operation [1:0] $end
$var wire 1 E3 Result $end
$var wire 1 F3 a $end
$var wire 1 G3 b $end
$var wire 2 H3 mux0inputs [1:0] $end
$var wire 2 I3 mux1inputs [1:0] $end
$var wire 4 J3 mux2inputs [3:0] $end
$var wire 1 K3 w1 $end
$var wire 1 L3 w2 $end
$scope module P0 $end
$var wire 2 M3 inputLines [1:0] $end
$var wire 1 K3 outputLine $end
$var wire 1 ?3 selectLine $end
$var wire 1 N3 w1 $end
$var wire 1 O3 w2 $end
$var wire 1 P3 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 Q3 inputLines [1:0] $end
$var wire 1 L3 outputLine $end
$var wire 1 @3 selectLine $end
$var wire 1 R3 w1 $end
$var wire 1 S3 w2 $end
$var wire 1 T3 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 K3 a $end
$var wire 1 L3 b $end
$var wire 1 A3 cin $end
$var wire 1 B3 cout $end
$var wire 1 U3 sum $end
$var wire 1 V3 w1 $end
$var wire 1 W3 w2 $end
$var wire 1 X3 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 Y3 inputLines [3:0] $end
$var wire 1 E3 outputLine $end
$var wire 2 Z3 selectLines [1:0] $end
$var wire 2 [3 w [1:0] $end
$scope module M0 $end
$var wire 2 \3 inputLines [1:0] $end
$var wire 1 ]3 outputLine $end
$var wire 1 ^3 selectLine $end
$var wire 1 _3 w1 $end
$var wire 1 `3 w2 $end
$var wire 1 a3 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 b3 inputLines [1:0] $end
$var wire 1 c3 outputLine $end
$var wire 1 d3 selectLine $end
$var wire 1 e3 w1 $end
$var wire 1 f3 w2 $end
$var wire 1 g3 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 h3 inputLines [1:0] $end
$var wire 1 E3 outputLine $end
$var wire 1 i3 selectLine $end
$var wire 1 j3 w1 $end
$var wire 1 k3 w2 $end
$var wire 1 l3 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A38 $end
$var wire 1 m3 Ainvert $end
$var wire 1 n3 Binvert $end
$var wire 1 o3 CarryIn $end
$var wire 1 p3 CarryOut $end
$var wire 1 q3 Less $end
$var wire 2 r3 Operation [1:0] $end
$var wire 1 s3 Result $end
$var wire 1 t3 a $end
$var wire 1 u3 b $end
$var wire 2 v3 mux0inputs [1:0] $end
$var wire 2 w3 mux1inputs [1:0] $end
$var wire 4 x3 mux2inputs [3:0] $end
$var wire 1 y3 w1 $end
$var wire 1 z3 w2 $end
$scope module P0 $end
$var wire 2 {3 inputLines [1:0] $end
$var wire 1 y3 outputLine $end
$var wire 1 m3 selectLine $end
$var wire 1 |3 w1 $end
$var wire 1 }3 w2 $end
$var wire 1 ~3 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 !4 inputLines [1:0] $end
$var wire 1 z3 outputLine $end
$var wire 1 n3 selectLine $end
$var wire 1 "4 w1 $end
$var wire 1 #4 w2 $end
$var wire 1 $4 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 y3 a $end
$var wire 1 z3 b $end
$var wire 1 o3 cin $end
$var wire 1 p3 cout $end
$var wire 1 %4 sum $end
$var wire 1 &4 w1 $end
$var wire 1 '4 w2 $end
$var wire 1 (4 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 )4 inputLines [3:0] $end
$var wire 1 s3 outputLine $end
$var wire 2 *4 selectLines [1:0] $end
$var wire 2 +4 w [1:0] $end
$scope module M0 $end
$var wire 2 ,4 inputLines [1:0] $end
$var wire 1 -4 outputLine $end
$var wire 1 .4 selectLine $end
$var wire 1 /4 w1 $end
$var wire 1 04 w2 $end
$var wire 1 14 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 24 inputLines [1:0] $end
$var wire 1 34 outputLine $end
$var wire 1 44 selectLine $end
$var wire 1 54 w1 $end
$var wire 1 64 w2 $end
$var wire 1 74 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 84 inputLines [1:0] $end
$var wire 1 s3 outputLine $end
$var wire 1 94 selectLine $end
$var wire 1 :4 w1 $end
$var wire 1 ;4 w2 $end
$var wire 1 <4 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A39 $end
$var wire 1 =4 Ainvert $end
$var wire 1 >4 Binvert $end
$var wire 1 ?4 CarryIn $end
$var wire 1 @4 CarryOut $end
$var wire 1 A4 Less $end
$var wire 2 B4 Operation [1:0] $end
$var wire 1 C4 Result $end
$var wire 1 D4 a $end
$var wire 1 E4 b $end
$var wire 2 F4 mux0inputs [1:0] $end
$var wire 2 G4 mux1inputs [1:0] $end
$var wire 4 H4 mux2inputs [3:0] $end
$var wire 1 I4 w1 $end
$var wire 1 J4 w2 $end
$scope module P0 $end
$var wire 2 K4 inputLines [1:0] $end
$var wire 1 I4 outputLine $end
$var wire 1 =4 selectLine $end
$var wire 1 L4 w1 $end
$var wire 1 M4 w2 $end
$var wire 1 N4 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 O4 inputLines [1:0] $end
$var wire 1 J4 outputLine $end
$var wire 1 >4 selectLine $end
$var wire 1 P4 w1 $end
$var wire 1 Q4 w2 $end
$var wire 1 R4 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 I4 a $end
$var wire 1 J4 b $end
$var wire 1 ?4 cin $end
$var wire 1 @4 cout $end
$var wire 1 S4 sum $end
$var wire 1 T4 w1 $end
$var wire 1 U4 w2 $end
$var wire 1 V4 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 W4 inputLines [3:0] $end
$var wire 1 C4 outputLine $end
$var wire 2 X4 selectLines [1:0] $end
$var wire 2 Y4 w [1:0] $end
$scope module M0 $end
$var wire 2 Z4 inputLines [1:0] $end
$var wire 1 [4 outputLine $end
$var wire 1 \4 selectLine $end
$var wire 1 ]4 w1 $end
$var wire 1 ^4 w2 $end
$var wire 1 _4 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 `4 inputLines [1:0] $end
$var wire 1 a4 outputLine $end
$var wire 1 b4 selectLine $end
$var wire 1 c4 w1 $end
$var wire 1 d4 w2 $end
$var wire 1 e4 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 f4 inputLines [1:0] $end
$var wire 1 C4 outputLine $end
$var wire 1 g4 selectLine $end
$var wire 1 h4 w1 $end
$var wire 1 i4 w2 $end
$var wire 1 j4 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A40 $end
$var wire 1 k4 Ainvert $end
$var wire 1 l4 Binvert $end
$var wire 1 m4 CarryIn $end
$var wire 1 n4 CarryOut $end
$var wire 1 o4 Less $end
$var wire 2 p4 Operation [1:0] $end
$var wire 1 q4 Result $end
$var wire 1 r4 a $end
$var wire 1 s4 b $end
$var wire 2 t4 mux0inputs [1:0] $end
$var wire 2 u4 mux1inputs [1:0] $end
$var wire 4 v4 mux2inputs [3:0] $end
$var wire 1 w4 w1 $end
$var wire 1 x4 w2 $end
$scope module P0 $end
$var wire 2 y4 inputLines [1:0] $end
$var wire 1 w4 outputLine $end
$var wire 1 k4 selectLine $end
$var wire 1 z4 w1 $end
$var wire 1 {4 w2 $end
$var wire 1 |4 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 }4 inputLines [1:0] $end
$var wire 1 x4 outputLine $end
$var wire 1 l4 selectLine $end
$var wire 1 ~4 w1 $end
$var wire 1 !5 w2 $end
$var wire 1 "5 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 w4 a $end
$var wire 1 x4 b $end
$var wire 1 m4 cin $end
$var wire 1 n4 cout $end
$var wire 1 #5 sum $end
$var wire 1 $5 w1 $end
$var wire 1 %5 w2 $end
$var wire 1 &5 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 '5 inputLines [3:0] $end
$var wire 1 q4 outputLine $end
$var wire 2 (5 selectLines [1:0] $end
$var wire 2 )5 w [1:0] $end
$scope module M0 $end
$var wire 2 *5 inputLines [1:0] $end
$var wire 1 +5 outputLine $end
$var wire 1 ,5 selectLine $end
$var wire 1 -5 w1 $end
$var wire 1 .5 w2 $end
$var wire 1 /5 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 05 inputLines [1:0] $end
$var wire 1 15 outputLine $end
$var wire 1 25 selectLine $end
$var wire 1 35 w1 $end
$var wire 1 45 w2 $end
$var wire 1 55 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 65 inputLines [1:0] $end
$var wire 1 q4 outputLine $end
$var wire 1 75 selectLine $end
$var wire 1 85 w1 $end
$var wire 1 95 w2 $end
$var wire 1 :5 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A41 $end
$var wire 1 ;5 Ainvert $end
$var wire 1 <5 Binvert $end
$var wire 1 =5 CarryIn $end
$var wire 1 >5 CarryOut $end
$var wire 1 ?5 Less $end
$var wire 2 @5 Operation [1:0] $end
$var wire 1 A5 Result $end
$var wire 1 B5 a $end
$var wire 1 C5 b $end
$var wire 2 D5 mux0inputs [1:0] $end
$var wire 2 E5 mux1inputs [1:0] $end
$var wire 4 F5 mux2inputs [3:0] $end
$var wire 1 G5 w1 $end
$var wire 1 H5 w2 $end
$scope module P0 $end
$var wire 2 I5 inputLines [1:0] $end
$var wire 1 G5 outputLine $end
$var wire 1 ;5 selectLine $end
$var wire 1 J5 w1 $end
$var wire 1 K5 w2 $end
$var wire 1 L5 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 M5 inputLines [1:0] $end
$var wire 1 H5 outputLine $end
$var wire 1 <5 selectLine $end
$var wire 1 N5 w1 $end
$var wire 1 O5 w2 $end
$var wire 1 P5 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 G5 a $end
$var wire 1 H5 b $end
$var wire 1 =5 cin $end
$var wire 1 >5 cout $end
$var wire 1 Q5 sum $end
$var wire 1 R5 w1 $end
$var wire 1 S5 w2 $end
$var wire 1 T5 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 U5 inputLines [3:0] $end
$var wire 1 A5 outputLine $end
$var wire 2 V5 selectLines [1:0] $end
$var wire 2 W5 w [1:0] $end
$scope module M0 $end
$var wire 2 X5 inputLines [1:0] $end
$var wire 1 Y5 outputLine $end
$var wire 1 Z5 selectLine $end
$var wire 1 [5 w1 $end
$var wire 1 \5 w2 $end
$var wire 1 ]5 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 ^5 inputLines [1:0] $end
$var wire 1 _5 outputLine $end
$var wire 1 `5 selectLine $end
$var wire 1 a5 w1 $end
$var wire 1 b5 w2 $end
$var wire 1 c5 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 d5 inputLines [1:0] $end
$var wire 1 A5 outputLine $end
$var wire 1 e5 selectLine $end
$var wire 1 f5 w1 $end
$var wire 1 g5 w2 $end
$var wire 1 h5 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A42 $end
$var wire 1 i5 Ainvert $end
$var wire 1 j5 Binvert $end
$var wire 1 k5 CarryIn $end
$var wire 1 l5 CarryOut $end
$var wire 1 m5 Less $end
$var wire 2 n5 Operation [1:0] $end
$var wire 1 o5 Result $end
$var wire 1 p5 a $end
$var wire 1 q5 b $end
$var wire 2 r5 mux0inputs [1:0] $end
$var wire 2 s5 mux1inputs [1:0] $end
$var wire 4 t5 mux2inputs [3:0] $end
$var wire 1 u5 w1 $end
$var wire 1 v5 w2 $end
$scope module P0 $end
$var wire 2 w5 inputLines [1:0] $end
$var wire 1 u5 outputLine $end
$var wire 1 i5 selectLine $end
$var wire 1 x5 w1 $end
$var wire 1 y5 w2 $end
$var wire 1 z5 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 {5 inputLines [1:0] $end
$var wire 1 v5 outputLine $end
$var wire 1 j5 selectLine $end
$var wire 1 |5 w1 $end
$var wire 1 }5 w2 $end
$var wire 1 ~5 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 u5 a $end
$var wire 1 v5 b $end
$var wire 1 k5 cin $end
$var wire 1 l5 cout $end
$var wire 1 !6 sum $end
$var wire 1 "6 w1 $end
$var wire 1 #6 w2 $end
$var wire 1 $6 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 %6 inputLines [3:0] $end
$var wire 1 o5 outputLine $end
$var wire 2 &6 selectLines [1:0] $end
$var wire 2 '6 w [1:0] $end
$scope module M0 $end
$var wire 2 (6 inputLines [1:0] $end
$var wire 1 )6 outputLine $end
$var wire 1 *6 selectLine $end
$var wire 1 +6 w1 $end
$var wire 1 ,6 w2 $end
$var wire 1 -6 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 .6 inputLines [1:0] $end
$var wire 1 /6 outputLine $end
$var wire 1 06 selectLine $end
$var wire 1 16 w1 $end
$var wire 1 26 w2 $end
$var wire 1 36 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 46 inputLines [1:0] $end
$var wire 1 o5 outputLine $end
$var wire 1 56 selectLine $end
$var wire 1 66 w1 $end
$var wire 1 76 w2 $end
$var wire 1 86 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A43 $end
$var wire 1 96 Ainvert $end
$var wire 1 :6 Binvert $end
$var wire 1 ;6 CarryIn $end
$var wire 1 <6 CarryOut $end
$var wire 1 =6 Less $end
$var wire 2 >6 Operation [1:0] $end
$var wire 1 ?6 Result $end
$var wire 1 @6 a $end
$var wire 1 A6 b $end
$var wire 2 B6 mux0inputs [1:0] $end
$var wire 2 C6 mux1inputs [1:0] $end
$var wire 4 D6 mux2inputs [3:0] $end
$var wire 1 E6 w1 $end
$var wire 1 F6 w2 $end
$scope module P0 $end
$var wire 2 G6 inputLines [1:0] $end
$var wire 1 E6 outputLine $end
$var wire 1 96 selectLine $end
$var wire 1 H6 w1 $end
$var wire 1 I6 w2 $end
$var wire 1 J6 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 K6 inputLines [1:0] $end
$var wire 1 F6 outputLine $end
$var wire 1 :6 selectLine $end
$var wire 1 L6 w1 $end
$var wire 1 M6 w2 $end
$var wire 1 N6 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 E6 a $end
$var wire 1 F6 b $end
$var wire 1 ;6 cin $end
$var wire 1 <6 cout $end
$var wire 1 O6 sum $end
$var wire 1 P6 w1 $end
$var wire 1 Q6 w2 $end
$var wire 1 R6 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 S6 inputLines [3:0] $end
$var wire 1 ?6 outputLine $end
$var wire 2 T6 selectLines [1:0] $end
$var wire 2 U6 w [1:0] $end
$scope module M0 $end
$var wire 2 V6 inputLines [1:0] $end
$var wire 1 W6 outputLine $end
$var wire 1 X6 selectLine $end
$var wire 1 Y6 w1 $end
$var wire 1 Z6 w2 $end
$var wire 1 [6 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 \6 inputLines [1:0] $end
$var wire 1 ]6 outputLine $end
$var wire 1 ^6 selectLine $end
$var wire 1 _6 w1 $end
$var wire 1 `6 w2 $end
$var wire 1 a6 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 b6 inputLines [1:0] $end
$var wire 1 ?6 outputLine $end
$var wire 1 c6 selectLine $end
$var wire 1 d6 w1 $end
$var wire 1 e6 w2 $end
$var wire 1 f6 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A44 $end
$var wire 1 g6 Ainvert $end
$var wire 1 h6 Binvert $end
$var wire 1 i6 CarryIn $end
$var wire 1 j6 CarryOut $end
$var wire 1 k6 Less $end
$var wire 2 l6 Operation [1:0] $end
$var wire 1 m6 Result $end
$var wire 1 n6 a $end
$var wire 1 o6 b $end
$var wire 2 p6 mux0inputs [1:0] $end
$var wire 2 q6 mux1inputs [1:0] $end
$var wire 4 r6 mux2inputs [3:0] $end
$var wire 1 s6 w1 $end
$var wire 1 t6 w2 $end
$scope module P0 $end
$var wire 2 u6 inputLines [1:0] $end
$var wire 1 s6 outputLine $end
$var wire 1 g6 selectLine $end
$var wire 1 v6 w1 $end
$var wire 1 w6 w2 $end
$var wire 1 x6 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 y6 inputLines [1:0] $end
$var wire 1 t6 outputLine $end
$var wire 1 h6 selectLine $end
$var wire 1 z6 w1 $end
$var wire 1 {6 w2 $end
$var wire 1 |6 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 s6 a $end
$var wire 1 t6 b $end
$var wire 1 i6 cin $end
$var wire 1 j6 cout $end
$var wire 1 }6 sum $end
$var wire 1 ~6 w1 $end
$var wire 1 !7 w2 $end
$var wire 1 "7 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 #7 inputLines [3:0] $end
$var wire 1 m6 outputLine $end
$var wire 2 $7 selectLines [1:0] $end
$var wire 2 %7 w [1:0] $end
$scope module M0 $end
$var wire 2 &7 inputLines [1:0] $end
$var wire 1 '7 outputLine $end
$var wire 1 (7 selectLine $end
$var wire 1 )7 w1 $end
$var wire 1 *7 w2 $end
$var wire 1 +7 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 ,7 inputLines [1:0] $end
$var wire 1 -7 outputLine $end
$var wire 1 .7 selectLine $end
$var wire 1 /7 w1 $end
$var wire 1 07 w2 $end
$var wire 1 17 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 27 inputLines [1:0] $end
$var wire 1 m6 outputLine $end
$var wire 1 37 selectLine $end
$var wire 1 47 w1 $end
$var wire 1 57 w2 $end
$var wire 1 67 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A45 $end
$var wire 1 77 Ainvert $end
$var wire 1 87 Binvert $end
$var wire 1 97 CarryIn $end
$var wire 1 :7 CarryOut $end
$var wire 1 ;7 Less $end
$var wire 2 <7 Operation [1:0] $end
$var wire 1 =7 Result $end
$var wire 1 >7 a $end
$var wire 1 ?7 b $end
$var wire 2 @7 mux0inputs [1:0] $end
$var wire 2 A7 mux1inputs [1:0] $end
$var wire 4 B7 mux2inputs [3:0] $end
$var wire 1 C7 w1 $end
$var wire 1 D7 w2 $end
$scope module P0 $end
$var wire 2 E7 inputLines [1:0] $end
$var wire 1 C7 outputLine $end
$var wire 1 77 selectLine $end
$var wire 1 F7 w1 $end
$var wire 1 G7 w2 $end
$var wire 1 H7 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 I7 inputLines [1:0] $end
$var wire 1 D7 outputLine $end
$var wire 1 87 selectLine $end
$var wire 1 J7 w1 $end
$var wire 1 K7 w2 $end
$var wire 1 L7 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 C7 a $end
$var wire 1 D7 b $end
$var wire 1 97 cin $end
$var wire 1 :7 cout $end
$var wire 1 M7 sum $end
$var wire 1 N7 w1 $end
$var wire 1 O7 w2 $end
$var wire 1 P7 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 Q7 inputLines [3:0] $end
$var wire 1 =7 outputLine $end
$var wire 2 R7 selectLines [1:0] $end
$var wire 2 S7 w [1:0] $end
$scope module M0 $end
$var wire 2 T7 inputLines [1:0] $end
$var wire 1 U7 outputLine $end
$var wire 1 V7 selectLine $end
$var wire 1 W7 w1 $end
$var wire 1 X7 w2 $end
$var wire 1 Y7 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 Z7 inputLines [1:0] $end
$var wire 1 [7 outputLine $end
$var wire 1 \7 selectLine $end
$var wire 1 ]7 w1 $end
$var wire 1 ^7 w2 $end
$var wire 1 _7 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 `7 inputLines [1:0] $end
$var wire 1 =7 outputLine $end
$var wire 1 a7 selectLine $end
$var wire 1 b7 w1 $end
$var wire 1 c7 w2 $end
$var wire 1 d7 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A46 $end
$var wire 1 e7 Ainvert $end
$var wire 1 f7 Binvert $end
$var wire 1 g7 CarryIn $end
$var wire 1 h7 CarryOut $end
$var wire 1 i7 Less $end
$var wire 2 j7 Operation [1:0] $end
$var wire 1 k7 Result $end
$var wire 1 l7 a $end
$var wire 1 m7 b $end
$var wire 2 n7 mux0inputs [1:0] $end
$var wire 2 o7 mux1inputs [1:0] $end
$var wire 4 p7 mux2inputs [3:0] $end
$var wire 1 q7 w1 $end
$var wire 1 r7 w2 $end
$scope module P0 $end
$var wire 2 s7 inputLines [1:0] $end
$var wire 1 q7 outputLine $end
$var wire 1 e7 selectLine $end
$var wire 1 t7 w1 $end
$var wire 1 u7 w2 $end
$var wire 1 v7 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 w7 inputLines [1:0] $end
$var wire 1 r7 outputLine $end
$var wire 1 f7 selectLine $end
$var wire 1 x7 w1 $end
$var wire 1 y7 w2 $end
$var wire 1 z7 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 q7 a $end
$var wire 1 r7 b $end
$var wire 1 g7 cin $end
$var wire 1 h7 cout $end
$var wire 1 {7 sum $end
$var wire 1 |7 w1 $end
$var wire 1 }7 w2 $end
$var wire 1 ~7 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 !8 inputLines [3:0] $end
$var wire 1 k7 outputLine $end
$var wire 2 "8 selectLines [1:0] $end
$var wire 2 #8 w [1:0] $end
$scope module M0 $end
$var wire 2 $8 inputLines [1:0] $end
$var wire 1 %8 outputLine $end
$var wire 1 &8 selectLine $end
$var wire 1 '8 w1 $end
$var wire 1 (8 w2 $end
$var wire 1 )8 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 *8 inputLines [1:0] $end
$var wire 1 +8 outputLine $end
$var wire 1 ,8 selectLine $end
$var wire 1 -8 w1 $end
$var wire 1 .8 w2 $end
$var wire 1 /8 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 08 inputLines [1:0] $end
$var wire 1 k7 outputLine $end
$var wire 1 18 selectLine $end
$var wire 1 28 w1 $end
$var wire 1 38 w2 $end
$var wire 1 48 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A47 $end
$var wire 1 58 Ainvert $end
$var wire 1 68 Binvert $end
$var wire 1 78 CarryIn $end
$var wire 1 88 CarryOut $end
$var wire 1 98 Less $end
$var wire 2 :8 Operation [1:0] $end
$var wire 1 ;8 Result $end
$var wire 1 <8 a $end
$var wire 1 =8 b $end
$var wire 2 >8 mux0inputs [1:0] $end
$var wire 2 ?8 mux1inputs [1:0] $end
$var wire 4 @8 mux2inputs [3:0] $end
$var wire 1 A8 w1 $end
$var wire 1 B8 w2 $end
$scope module P0 $end
$var wire 2 C8 inputLines [1:0] $end
$var wire 1 A8 outputLine $end
$var wire 1 58 selectLine $end
$var wire 1 D8 w1 $end
$var wire 1 E8 w2 $end
$var wire 1 F8 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 G8 inputLines [1:0] $end
$var wire 1 B8 outputLine $end
$var wire 1 68 selectLine $end
$var wire 1 H8 w1 $end
$var wire 1 I8 w2 $end
$var wire 1 J8 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 A8 a $end
$var wire 1 B8 b $end
$var wire 1 78 cin $end
$var wire 1 88 cout $end
$var wire 1 K8 sum $end
$var wire 1 L8 w1 $end
$var wire 1 M8 w2 $end
$var wire 1 N8 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 O8 inputLines [3:0] $end
$var wire 1 ;8 outputLine $end
$var wire 2 P8 selectLines [1:0] $end
$var wire 2 Q8 w [1:0] $end
$scope module M0 $end
$var wire 2 R8 inputLines [1:0] $end
$var wire 1 S8 outputLine $end
$var wire 1 T8 selectLine $end
$var wire 1 U8 w1 $end
$var wire 1 V8 w2 $end
$var wire 1 W8 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 X8 inputLines [1:0] $end
$var wire 1 Y8 outputLine $end
$var wire 1 Z8 selectLine $end
$var wire 1 [8 w1 $end
$var wire 1 \8 w2 $end
$var wire 1 ]8 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 ^8 inputLines [1:0] $end
$var wire 1 ;8 outputLine $end
$var wire 1 _8 selectLine $end
$var wire 1 `8 w1 $end
$var wire 1 a8 w2 $end
$var wire 1 b8 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A48 $end
$var wire 1 c8 Ainvert $end
$var wire 1 d8 Binvert $end
$var wire 1 e8 CarryIn $end
$var wire 1 f8 CarryOut $end
$var wire 1 g8 Less $end
$var wire 2 h8 Operation [1:0] $end
$var wire 1 i8 Result $end
$var wire 1 j8 a $end
$var wire 1 k8 b $end
$var wire 2 l8 mux0inputs [1:0] $end
$var wire 2 m8 mux1inputs [1:0] $end
$var wire 4 n8 mux2inputs [3:0] $end
$var wire 1 o8 w1 $end
$var wire 1 p8 w2 $end
$scope module P0 $end
$var wire 2 q8 inputLines [1:0] $end
$var wire 1 o8 outputLine $end
$var wire 1 c8 selectLine $end
$var wire 1 r8 w1 $end
$var wire 1 s8 w2 $end
$var wire 1 t8 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 u8 inputLines [1:0] $end
$var wire 1 p8 outputLine $end
$var wire 1 d8 selectLine $end
$var wire 1 v8 w1 $end
$var wire 1 w8 w2 $end
$var wire 1 x8 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 o8 a $end
$var wire 1 p8 b $end
$var wire 1 e8 cin $end
$var wire 1 f8 cout $end
$var wire 1 y8 sum $end
$var wire 1 z8 w1 $end
$var wire 1 {8 w2 $end
$var wire 1 |8 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 }8 inputLines [3:0] $end
$var wire 1 i8 outputLine $end
$var wire 2 ~8 selectLines [1:0] $end
$var wire 2 !9 w [1:0] $end
$scope module M0 $end
$var wire 2 "9 inputLines [1:0] $end
$var wire 1 #9 outputLine $end
$var wire 1 $9 selectLine $end
$var wire 1 %9 w1 $end
$var wire 1 &9 w2 $end
$var wire 1 '9 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 (9 inputLines [1:0] $end
$var wire 1 )9 outputLine $end
$var wire 1 *9 selectLine $end
$var wire 1 +9 w1 $end
$var wire 1 ,9 w2 $end
$var wire 1 -9 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 .9 inputLines [1:0] $end
$var wire 1 i8 outputLine $end
$var wire 1 /9 selectLine $end
$var wire 1 09 w1 $end
$var wire 1 19 w2 $end
$var wire 1 29 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A49 $end
$var wire 1 39 Ainvert $end
$var wire 1 49 Binvert $end
$var wire 1 59 CarryIn $end
$var wire 1 69 CarryOut $end
$var wire 1 79 Less $end
$var wire 2 89 Operation [1:0] $end
$var wire 1 99 Result $end
$var wire 1 :9 a $end
$var wire 1 ;9 b $end
$var wire 2 <9 mux0inputs [1:0] $end
$var wire 2 =9 mux1inputs [1:0] $end
$var wire 4 >9 mux2inputs [3:0] $end
$var wire 1 ?9 w1 $end
$var wire 1 @9 w2 $end
$scope module P0 $end
$var wire 2 A9 inputLines [1:0] $end
$var wire 1 ?9 outputLine $end
$var wire 1 39 selectLine $end
$var wire 1 B9 w1 $end
$var wire 1 C9 w2 $end
$var wire 1 D9 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 E9 inputLines [1:0] $end
$var wire 1 @9 outputLine $end
$var wire 1 49 selectLine $end
$var wire 1 F9 w1 $end
$var wire 1 G9 w2 $end
$var wire 1 H9 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 ?9 a $end
$var wire 1 @9 b $end
$var wire 1 59 cin $end
$var wire 1 69 cout $end
$var wire 1 I9 sum $end
$var wire 1 J9 w1 $end
$var wire 1 K9 w2 $end
$var wire 1 L9 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 M9 inputLines [3:0] $end
$var wire 1 99 outputLine $end
$var wire 2 N9 selectLines [1:0] $end
$var wire 2 O9 w [1:0] $end
$scope module M0 $end
$var wire 2 P9 inputLines [1:0] $end
$var wire 1 Q9 outputLine $end
$var wire 1 R9 selectLine $end
$var wire 1 S9 w1 $end
$var wire 1 T9 w2 $end
$var wire 1 U9 w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 V9 inputLines [1:0] $end
$var wire 1 W9 outputLine $end
$var wire 1 X9 selectLine $end
$var wire 1 Y9 w1 $end
$var wire 1 Z9 w2 $end
$var wire 1 [9 w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 \9 inputLines [1:0] $end
$var wire 1 99 outputLine $end
$var wire 1 ]9 selectLine $end
$var wire 1 ^9 w1 $end
$var wire 1 _9 w2 $end
$var wire 1 `9 w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A50 $end
$var wire 1 a9 Ainvert $end
$var wire 1 b9 Binvert $end
$var wire 1 c9 CarryIn $end
$var wire 1 d9 CarryOut $end
$var wire 1 e9 Less $end
$var wire 2 f9 Operation [1:0] $end
$var wire 1 g9 Result $end
$var wire 1 h9 a $end
$var wire 1 i9 b $end
$var wire 2 j9 mux0inputs [1:0] $end
$var wire 2 k9 mux1inputs [1:0] $end
$var wire 4 l9 mux2inputs [3:0] $end
$var wire 1 m9 w1 $end
$var wire 1 n9 w2 $end
$scope module P0 $end
$var wire 2 o9 inputLines [1:0] $end
$var wire 1 m9 outputLine $end
$var wire 1 a9 selectLine $end
$var wire 1 p9 w1 $end
$var wire 1 q9 w2 $end
$var wire 1 r9 w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 s9 inputLines [1:0] $end
$var wire 1 n9 outputLine $end
$var wire 1 b9 selectLine $end
$var wire 1 t9 w1 $end
$var wire 1 u9 w2 $end
$var wire 1 v9 w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 m9 a $end
$var wire 1 n9 b $end
$var wire 1 c9 cin $end
$var wire 1 d9 cout $end
$var wire 1 w9 sum $end
$var wire 1 x9 w1 $end
$var wire 1 y9 w2 $end
$var wire 1 z9 w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 {9 inputLines [3:0] $end
$var wire 1 g9 outputLine $end
$var wire 2 |9 selectLines [1:0] $end
$var wire 2 }9 w [1:0] $end
$scope module M0 $end
$var wire 2 ~9 inputLines [1:0] $end
$var wire 1 !: outputLine $end
$var wire 1 ": selectLine $end
$var wire 1 #: w1 $end
$var wire 1 $: w2 $end
$var wire 1 %: w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 &: inputLines [1:0] $end
$var wire 1 ': outputLine $end
$var wire 1 (: selectLine $end
$var wire 1 ): w1 $end
$var wire 1 *: w2 $end
$var wire 1 +: w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 ,: inputLines [1:0] $end
$var wire 1 g9 outputLine $end
$var wire 1 -: selectLine $end
$var wire 1 .: w1 $end
$var wire 1 /: w2 $end
$var wire 1 0: w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A51 $end
$var wire 1 1: Ainvert $end
$var wire 1 2: Binvert $end
$var wire 1 3: CarryIn $end
$var wire 1 4: CarryOut $end
$var wire 1 5: Less $end
$var wire 2 6: Operation [1:0] $end
$var wire 1 7: Result $end
$var wire 1 8: a $end
$var wire 1 9: b $end
$var wire 2 :: mux0inputs [1:0] $end
$var wire 2 ;: mux1inputs [1:0] $end
$var wire 4 <: mux2inputs [3:0] $end
$var wire 1 =: w1 $end
$var wire 1 >: w2 $end
$scope module P0 $end
$var wire 2 ?: inputLines [1:0] $end
$var wire 1 =: outputLine $end
$var wire 1 1: selectLine $end
$var wire 1 @: w1 $end
$var wire 1 A: w2 $end
$var wire 1 B: w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 C: inputLines [1:0] $end
$var wire 1 >: outputLine $end
$var wire 1 2: selectLine $end
$var wire 1 D: w1 $end
$var wire 1 E: w2 $end
$var wire 1 F: w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 =: a $end
$var wire 1 >: b $end
$var wire 1 3: cin $end
$var wire 1 4: cout $end
$var wire 1 G: sum $end
$var wire 1 H: w1 $end
$var wire 1 I: w2 $end
$var wire 1 J: w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 K: inputLines [3:0] $end
$var wire 1 7: outputLine $end
$var wire 2 L: selectLines [1:0] $end
$var wire 2 M: w [1:0] $end
$scope module M0 $end
$var wire 2 N: inputLines [1:0] $end
$var wire 1 O: outputLine $end
$var wire 1 P: selectLine $end
$var wire 1 Q: w1 $end
$var wire 1 R: w2 $end
$var wire 1 S: w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 T: inputLines [1:0] $end
$var wire 1 U: outputLine $end
$var wire 1 V: selectLine $end
$var wire 1 W: w1 $end
$var wire 1 X: w2 $end
$var wire 1 Y: w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 Z: inputLines [1:0] $end
$var wire 1 7: outputLine $end
$var wire 1 [: selectLine $end
$var wire 1 \: w1 $end
$var wire 1 ]: w2 $end
$var wire 1 ^: w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A52 $end
$var wire 1 _: Ainvert $end
$var wire 1 `: Binvert $end
$var wire 1 a: CarryIn $end
$var wire 1 b: CarryOut $end
$var wire 1 c: Less $end
$var wire 2 d: Operation [1:0] $end
$var wire 1 e: Result $end
$var wire 1 f: a $end
$var wire 1 g: b $end
$var wire 2 h: mux0inputs [1:0] $end
$var wire 2 i: mux1inputs [1:0] $end
$var wire 4 j: mux2inputs [3:0] $end
$var wire 1 k: w1 $end
$var wire 1 l: w2 $end
$scope module P0 $end
$var wire 2 m: inputLines [1:0] $end
$var wire 1 k: outputLine $end
$var wire 1 _: selectLine $end
$var wire 1 n: w1 $end
$var wire 1 o: w2 $end
$var wire 1 p: w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 q: inputLines [1:0] $end
$var wire 1 l: outputLine $end
$var wire 1 `: selectLine $end
$var wire 1 r: w1 $end
$var wire 1 s: w2 $end
$var wire 1 t: w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 k: a $end
$var wire 1 l: b $end
$var wire 1 a: cin $end
$var wire 1 b: cout $end
$var wire 1 u: sum $end
$var wire 1 v: w1 $end
$var wire 1 w: w2 $end
$var wire 1 x: w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 y: inputLines [3:0] $end
$var wire 1 e: outputLine $end
$var wire 2 z: selectLines [1:0] $end
$var wire 2 {: w [1:0] $end
$scope module M0 $end
$var wire 2 |: inputLines [1:0] $end
$var wire 1 }: outputLine $end
$var wire 1 ~: selectLine $end
$var wire 1 !; w1 $end
$var wire 1 "; w2 $end
$var wire 1 #; w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 $; inputLines [1:0] $end
$var wire 1 %; outputLine $end
$var wire 1 &; selectLine $end
$var wire 1 '; w1 $end
$var wire 1 (; w2 $end
$var wire 1 ); w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 *; inputLines [1:0] $end
$var wire 1 e: outputLine $end
$var wire 1 +; selectLine $end
$var wire 1 ,; w1 $end
$var wire 1 -; w2 $end
$var wire 1 .; w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A53 $end
$var wire 1 /; Ainvert $end
$var wire 1 0; Binvert $end
$var wire 1 1; CarryIn $end
$var wire 1 2; CarryOut $end
$var wire 1 3; Less $end
$var wire 2 4; Operation [1:0] $end
$var wire 1 5; Result $end
$var wire 1 6; a $end
$var wire 1 7; b $end
$var wire 2 8; mux0inputs [1:0] $end
$var wire 2 9; mux1inputs [1:0] $end
$var wire 4 :; mux2inputs [3:0] $end
$var wire 1 ;; w1 $end
$var wire 1 <; w2 $end
$scope module P0 $end
$var wire 2 =; inputLines [1:0] $end
$var wire 1 ;; outputLine $end
$var wire 1 /; selectLine $end
$var wire 1 >; w1 $end
$var wire 1 ?; w2 $end
$var wire 1 @; w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 A; inputLines [1:0] $end
$var wire 1 <; outputLine $end
$var wire 1 0; selectLine $end
$var wire 1 B; w1 $end
$var wire 1 C; w2 $end
$var wire 1 D; w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 ;; a $end
$var wire 1 <; b $end
$var wire 1 1; cin $end
$var wire 1 2; cout $end
$var wire 1 E; sum $end
$var wire 1 F; w1 $end
$var wire 1 G; w2 $end
$var wire 1 H; w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 I; inputLines [3:0] $end
$var wire 1 5; outputLine $end
$var wire 2 J; selectLines [1:0] $end
$var wire 2 K; w [1:0] $end
$scope module M0 $end
$var wire 2 L; inputLines [1:0] $end
$var wire 1 M; outputLine $end
$var wire 1 N; selectLine $end
$var wire 1 O; w1 $end
$var wire 1 P; w2 $end
$var wire 1 Q; w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 R; inputLines [1:0] $end
$var wire 1 S; outputLine $end
$var wire 1 T; selectLine $end
$var wire 1 U; w1 $end
$var wire 1 V; w2 $end
$var wire 1 W; w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 X; inputLines [1:0] $end
$var wire 1 5; outputLine $end
$var wire 1 Y; selectLine $end
$var wire 1 Z; w1 $end
$var wire 1 [; w2 $end
$var wire 1 \; w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A54 $end
$var wire 1 ]; Ainvert $end
$var wire 1 ^; Binvert $end
$var wire 1 _; CarryIn $end
$var wire 1 `; CarryOut $end
$var wire 1 a; Less $end
$var wire 2 b; Operation [1:0] $end
$var wire 1 c; Result $end
$var wire 1 d; a $end
$var wire 1 e; b $end
$var wire 2 f; mux0inputs [1:0] $end
$var wire 2 g; mux1inputs [1:0] $end
$var wire 4 h; mux2inputs [3:0] $end
$var wire 1 i; w1 $end
$var wire 1 j; w2 $end
$scope module P0 $end
$var wire 2 k; inputLines [1:0] $end
$var wire 1 i; outputLine $end
$var wire 1 ]; selectLine $end
$var wire 1 l; w1 $end
$var wire 1 m; w2 $end
$var wire 1 n; w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 o; inputLines [1:0] $end
$var wire 1 j; outputLine $end
$var wire 1 ^; selectLine $end
$var wire 1 p; w1 $end
$var wire 1 q; w2 $end
$var wire 1 r; w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 i; a $end
$var wire 1 j; b $end
$var wire 1 _; cin $end
$var wire 1 `; cout $end
$var wire 1 s; sum $end
$var wire 1 t; w1 $end
$var wire 1 u; w2 $end
$var wire 1 v; w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 w; inputLines [3:0] $end
$var wire 1 c; outputLine $end
$var wire 2 x; selectLines [1:0] $end
$var wire 2 y; w [1:0] $end
$scope module M0 $end
$var wire 2 z; inputLines [1:0] $end
$var wire 1 {; outputLine $end
$var wire 1 |; selectLine $end
$var wire 1 }; w1 $end
$var wire 1 ~; w2 $end
$var wire 1 !< w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 "< inputLines [1:0] $end
$var wire 1 #< outputLine $end
$var wire 1 $< selectLine $end
$var wire 1 %< w1 $end
$var wire 1 &< w2 $end
$var wire 1 '< w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 (< inputLines [1:0] $end
$var wire 1 c; outputLine $end
$var wire 1 )< selectLine $end
$var wire 1 *< w1 $end
$var wire 1 +< w2 $end
$var wire 1 ,< w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A55 $end
$var wire 1 -< Ainvert $end
$var wire 1 .< Binvert $end
$var wire 1 /< CarryIn $end
$var wire 1 0< CarryOut $end
$var wire 1 1< Less $end
$var wire 2 2< Operation [1:0] $end
$var wire 1 3< Result $end
$var wire 1 4< a $end
$var wire 1 5< b $end
$var wire 2 6< mux0inputs [1:0] $end
$var wire 2 7< mux1inputs [1:0] $end
$var wire 4 8< mux2inputs [3:0] $end
$var wire 1 9< w1 $end
$var wire 1 :< w2 $end
$scope module P0 $end
$var wire 2 ;< inputLines [1:0] $end
$var wire 1 9< outputLine $end
$var wire 1 -< selectLine $end
$var wire 1 << w1 $end
$var wire 1 =< w2 $end
$var wire 1 >< w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 ?< inputLines [1:0] $end
$var wire 1 :< outputLine $end
$var wire 1 .< selectLine $end
$var wire 1 @< w1 $end
$var wire 1 A< w2 $end
$var wire 1 B< w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 9< a $end
$var wire 1 :< b $end
$var wire 1 /< cin $end
$var wire 1 0< cout $end
$var wire 1 C< sum $end
$var wire 1 D< w1 $end
$var wire 1 E< w2 $end
$var wire 1 F< w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 G< inputLines [3:0] $end
$var wire 1 3< outputLine $end
$var wire 2 H< selectLines [1:0] $end
$var wire 2 I< w [1:0] $end
$scope module M0 $end
$var wire 2 J< inputLines [1:0] $end
$var wire 1 K< outputLine $end
$var wire 1 L< selectLine $end
$var wire 1 M< w1 $end
$var wire 1 N< w2 $end
$var wire 1 O< w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 P< inputLines [1:0] $end
$var wire 1 Q< outputLine $end
$var wire 1 R< selectLine $end
$var wire 1 S< w1 $end
$var wire 1 T< w2 $end
$var wire 1 U< w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 V< inputLines [1:0] $end
$var wire 1 3< outputLine $end
$var wire 1 W< selectLine $end
$var wire 1 X< w1 $end
$var wire 1 Y< w2 $end
$var wire 1 Z< w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A56 $end
$var wire 1 [< Ainvert $end
$var wire 1 \< Binvert $end
$var wire 1 ]< CarryIn $end
$var wire 1 ^< CarryOut $end
$var wire 1 _< Less $end
$var wire 2 `< Operation [1:0] $end
$var wire 1 a< Result $end
$var wire 1 b< a $end
$var wire 1 c< b $end
$var wire 2 d< mux0inputs [1:0] $end
$var wire 2 e< mux1inputs [1:0] $end
$var wire 4 f< mux2inputs [3:0] $end
$var wire 1 g< w1 $end
$var wire 1 h< w2 $end
$scope module P0 $end
$var wire 2 i< inputLines [1:0] $end
$var wire 1 g< outputLine $end
$var wire 1 [< selectLine $end
$var wire 1 j< w1 $end
$var wire 1 k< w2 $end
$var wire 1 l< w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 m< inputLines [1:0] $end
$var wire 1 h< outputLine $end
$var wire 1 \< selectLine $end
$var wire 1 n< w1 $end
$var wire 1 o< w2 $end
$var wire 1 p< w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 g< a $end
$var wire 1 h< b $end
$var wire 1 ]< cin $end
$var wire 1 ^< cout $end
$var wire 1 q< sum $end
$var wire 1 r< w1 $end
$var wire 1 s< w2 $end
$var wire 1 t< w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 u< inputLines [3:0] $end
$var wire 1 a< outputLine $end
$var wire 2 v< selectLines [1:0] $end
$var wire 2 w< w [1:0] $end
$scope module M0 $end
$var wire 2 x< inputLines [1:0] $end
$var wire 1 y< outputLine $end
$var wire 1 z< selectLine $end
$var wire 1 {< w1 $end
$var wire 1 |< w2 $end
$var wire 1 }< w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 ~< inputLines [1:0] $end
$var wire 1 != outputLine $end
$var wire 1 "= selectLine $end
$var wire 1 #= w1 $end
$var wire 1 $= w2 $end
$var wire 1 %= w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 &= inputLines [1:0] $end
$var wire 1 a< outputLine $end
$var wire 1 '= selectLine $end
$var wire 1 (= w1 $end
$var wire 1 )= w2 $end
$var wire 1 *= w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A57 $end
$var wire 1 += Ainvert $end
$var wire 1 ,= Binvert $end
$var wire 1 -= CarryIn $end
$var wire 1 .= CarryOut $end
$var wire 1 /= Less $end
$var wire 2 0= Operation [1:0] $end
$var wire 1 1= Result $end
$var wire 1 2= a $end
$var wire 1 3= b $end
$var wire 2 4= mux0inputs [1:0] $end
$var wire 2 5= mux1inputs [1:0] $end
$var wire 4 6= mux2inputs [3:0] $end
$var wire 1 7= w1 $end
$var wire 1 8= w2 $end
$scope module P0 $end
$var wire 2 9= inputLines [1:0] $end
$var wire 1 7= outputLine $end
$var wire 1 += selectLine $end
$var wire 1 := w1 $end
$var wire 1 ;= w2 $end
$var wire 1 <= w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 == inputLines [1:0] $end
$var wire 1 8= outputLine $end
$var wire 1 ,= selectLine $end
$var wire 1 >= w1 $end
$var wire 1 ?= w2 $end
$var wire 1 @= w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 7= a $end
$var wire 1 8= b $end
$var wire 1 -= cin $end
$var wire 1 .= cout $end
$var wire 1 A= sum $end
$var wire 1 B= w1 $end
$var wire 1 C= w2 $end
$var wire 1 D= w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 E= inputLines [3:0] $end
$var wire 1 1= outputLine $end
$var wire 2 F= selectLines [1:0] $end
$var wire 2 G= w [1:0] $end
$scope module M0 $end
$var wire 2 H= inputLines [1:0] $end
$var wire 1 I= outputLine $end
$var wire 1 J= selectLine $end
$var wire 1 K= w1 $end
$var wire 1 L= w2 $end
$var wire 1 M= w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 N= inputLines [1:0] $end
$var wire 1 O= outputLine $end
$var wire 1 P= selectLine $end
$var wire 1 Q= w1 $end
$var wire 1 R= w2 $end
$var wire 1 S= w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 T= inputLines [1:0] $end
$var wire 1 1= outputLine $end
$var wire 1 U= selectLine $end
$var wire 1 V= w1 $end
$var wire 1 W= w2 $end
$var wire 1 X= w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A58 $end
$var wire 1 Y= Ainvert $end
$var wire 1 Z= Binvert $end
$var wire 1 [= CarryIn $end
$var wire 1 \= CarryOut $end
$var wire 1 ]= Less $end
$var wire 2 ^= Operation [1:0] $end
$var wire 1 _= Result $end
$var wire 1 `= a $end
$var wire 1 a= b $end
$var wire 2 b= mux0inputs [1:0] $end
$var wire 2 c= mux1inputs [1:0] $end
$var wire 4 d= mux2inputs [3:0] $end
$var wire 1 e= w1 $end
$var wire 1 f= w2 $end
$scope module P0 $end
$var wire 2 g= inputLines [1:0] $end
$var wire 1 e= outputLine $end
$var wire 1 Y= selectLine $end
$var wire 1 h= w1 $end
$var wire 1 i= w2 $end
$var wire 1 j= w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 k= inputLines [1:0] $end
$var wire 1 f= outputLine $end
$var wire 1 Z= selectLine $end
$var wire 1 l= w1 $end
$var wire 1 m= w2 $end
$var wire 1 n= w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 e= a $end
$var wire 1 f= b $end
$var wire 1 [= cin $end
$var wire 1 \= cout $end
$var wire 1 o= sum $end
$var wire 1 p= w1 $end
$var wire 1 q= w2 $end
$var wire 1 r= w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 s= inputLines [3:0] $end
$var wire 1 _= outputLine $end
$var wire 2 t= selectLines [1:0] $end
$var wire 2 u= w [1:0] $end
$scope module M0 $end
$var wire 2 v= inputLines [1:0] $end
$var wire 1 w= outputLine $end
$var wire 1 x= selectLine $end
$var wire 1 y= w1 $end
$var wire 1 z= w2 $end
$var wire 1 {= w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 |= inputLines [1:0] $end
$var wire 1 }= outputLine $end
$var wire 1 ~= selectLine $end
$var wire 1 !> w1 $end
$var wire 1 "> w2 $end
$var wire 1 #> w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 $> inputLines [1:0] $end
$var wire 1 _= outputLine $end
$var wire 1 %> selectLine $end
$var wire 1 &> w1 $end
$var wire 1 '> w2 $end
$var wire 1 (> w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A59 $end
$var wire 1 )> Ainvert $end
$var wire 1 *> Binvert $end
$var wire 1 +> CarryIn $end
$var wire 1 ,> CarryOut $end
$var wire 1 -> Less $end
$var wire 2 .> Operation [1:0] $end
$var wire 1 /> Result $end
$var wire 1 0> a $end
$var wire 1 1> b $end
$var wire 2 2> mux0inputs [1:0] $end
$var wire 2 3> mux1inputs [1:0] $end
$var wire 4 4> mux2inputs [3:0] $end
$var wire 1 5> w1 $end
$var wire 1 6> w2 $end
$scope module P0 $end
$var wire 2 7> inputLines [1:0] $end
$var wire 1 5> outputLine $end
$var wire 1 )> selectLine $end
$var wire 1 8> w1 $end
$var wire 1 9> w2 $end
$var wire 1 :> w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 ;> inputLines [1:0] $end
$var wire 1 6> outputLine $end
$var wire 1 *> selectLine $end
$var wire 1 <> w1 $end
$var wire 1 => w2 $end
$var wire 1 >> w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 5> a $end
$var wire 1 6> b $end
$var wire 1 +> cin $end
$var wire 1 ,> cout $end
$var wire 1 ?> sum $end
$var wire 1 @> w1 $end
$var wire 1 A> w2 $end
$var wire 1 B> w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 C> inputLines [3:0] $end
$var wire 1 /> outputLine $end
$var wire 2 D> selectLines [1:0] $end
$var wire 2 E> w [1:0] $end
$scope module M0 $end
$var wire 2 F> inputLines [1:0] $end
$var wire 1 G> outputLine $end
$var wire 1 H> selectLine $end
$var wire 1 I> w1 $end
$var wire 1 J> w2 $end
$var wire 1 K> w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 L> inputLines [1:0] $end
$var wire 1 M> outputLine $end
$var wire 1 N> selectLine $end
$var wire 1 O> w1 $end
$var wire 1 P> w2 $end
$var wire 1 Q> w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 R> inputLines [1:0] $end
$var wire 1 /> outputLine $end
$var wire 1 S> selectLine $end
$var wire 1 T> w1 $end
$var wire 1 U> w2 $end
$var wire 1 V> w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A60 $end
$var wire 1 W> Ainvert $end
$var wire 1 X> Binvert $end
$var wire 1 Y> CarryIn $end
$var wire 1 Z> CarryOut $end
$var wire 1 [> Less $end
$var wire 2 \> Operation [1:0] $end
$var wire 1 ]> Result $end
$var wire 1 ^> a $end
$var wire 1 _> b $end
$var wire 2 `> mux0inputs [1:0] $end
$var wire 2 a> mux1inputs [1:0] $end
$var wire 4 b> mux2inputs [3:0] $end
$var wire 1 c> w1 $end
$var wire 1 d> w2 $end
$scope module P0 $end
$var wire 2 e> inputLines [1:0] $end
$var wire 1 c> outputLine $end
$var wire 1 W> selectLine $end
$var wire 1 f> w1 $end
$var wire 1 g> w2 $end
$var wire 1 h> w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 i> inputLines [1:0] $end
$var wire 1 d> outputLine $end
$var wire 1 X> selectLine $end
$var wire 1 j> w1 $end
$var wire 1 k> w2 $end
$var wire 1 l> w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 c> a $end
$var wire 1 d> b $end
$var wire 1 Y> cin $end
$var wire 1 Z> cout $end
$var wire 1 m> sum $end
$var wire 1 n> w1 $end
$var wire 1 o> w2 $end
$var wire 1 p> w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 q> inputLines [3:0] $end
$var wire 1 ]> outputLine $end
$var wire 2 r> selectLines [1:0] $end
$var wire 2 s> w [1:0] $end
$scope module M0 $end
$var wire 2 t> inputLines [1:0] $end
$var wire 1 u> outputLine $end
$var wire 1 v> selectLine $end
$var wire 1 w> w1 $end
$var wire 1 x> w2 $end
$var wire 1 y> w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 z> inputLines [1:0] $end
$var wire 1 {> outputLine $end
$var wire 1 |> selectLine $end
$var wire 1 }> w1 $end
$var wire 1 ~> w2 $end
$var wire 1 !? w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 "? inputLines [1:0] $end
$var wire 1 ]> outputLine $end
$var wire 1 #? selectLine $end
$var wire 1 $? w1 $end
$var wire 1 %? w2 $end
$var wire 1 &? w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A61 $end
$var wire 1 '? Ainvert $end
$var wire 1 (? Binvert $end
$var wire 1 )? CarryIn $end
$var wire 1 *? CarryOut $end
$var wire 1 +? Less $end
$var wire 2 ,? Operation [1:0] $end
$var wire 1 -? Result $end
$var wire 1 .? a $end
$var wire 1 /? b $end
$var wire 2 0? mux0inputs [1:0] $end
$var wire 2 1? mux1inputs [1:0] $end
$var wire 4 2? mux2inputs [3:0] $end
$var wire 1 3? w1 $end
$var wire 1 4? w2 $end
$scope module P0 $end
$var wire 2 5? inputLines [1:0] $end
$var wire 1 3? outputLine $end
$var wire 1 '? selectLine $end
$var wire 1 6? w1 $end
$var wire 1 7? w2 $end
$var wire 1 8? w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 9? inputLines [1:0] $end
$var wire 1 4? outputLine $end
$var wire 1 (? selectLine $end
$var wire 1 :? w1 $end
$var wire 1 ;? w2 $end
$var wire 1 <? w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 3? a $end
$var wire 1 4? b $end
$var wire 1 )? cin $end
$var wire 1 *? cout $end
$var wire 1 =? sum $end
$var wire 1 >? w1 $end
$var wire 1 ?? w2 $end
$var wire 1 @? w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 A? inputLines [3:0] $end
$var wire 1 -? outputLine $end
$var wire 2 B? selectLines [1:0] $end
$var wire 2 C? w [1:0] $end
$scope module M0 $end
$var wire 2 D? inputLines [1:0] $end
$var wire 1 E? outputLine $end
$var wire 1 F? selectLine $end
$var wire 1 G? w1 $end
$var wire 1 H? w2 $end
$var wire 1 I? w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 J? inputLines [1:0] $end
$var wire 1 K? outputLine $end
$var wire 1 L? selectLine $end
$var wire 1 M? w1 $end
$var wire 1 N? w2 $end
$var wire 1 O? w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 P? inputLines [1:0] $end
$var wire 1 -? outputLine $end
$var wire 1 Q? selectLine $end
$var wire 1 R? w1 $end
$var wire 1 S? w2 $end
$var wire 1 T? w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A62 $end
$var wire 1 U? Ainvert $end
$var wire 1 V? Binvert $end
$var wire 1 W? CarryIn $end
$var wire 1 X? CarryOut $end
$var wire 1 Y? Less $end
$var wire 2 Z? Operation [1:0] $end
$var wire 1 [? Result $end
$var wire 1 \? a $end
$var wire 1 ]? b $end
$var wire 2 ^? mux0inputs [1:0] $end
$var wire 2 _? mux1inputs [1:0] $end
$var wire 4 `? mux2inputs [3:0] $end
$var wire 1 a? w1 $end
$var wire 1 b? w2 $end
$scope module P0 $end
$var wire 2 c? inputLines [1:0] $end
$var wire 1 a? outputLine $end
$var wire 1 U? selectLine $end
$var wire 1 d? w1 $end
$var wire 1 e? w2 $end
$var wire 1 f? w3 $end
$upscope $end
$scope module P1 $end
$var wire 2 g? inputLines [1:0] $end
$var wire 1 b? outputLine $end
$var wire 1 V? selectLine $end
$var wire 1 h? w1 $end
$var wire 1 i? w2 $end
$var wire 1 j? w3 $end
$upscope $end
$scope module P4 $end
$var wire 1 a? a $end
$var wire 1 b? b $end
$var wire 1 W? cin $end
$var wire 1 X? cout $end
$var wire 1 k? sum $end
$var wire 1 l? w1 $end
$var wire 1 m? w2 $end
$var wire 1 n? w3 $end
$upscope $end
$scope module P5 $end
$var wire 4 o? inputLines [3:0] $end
$var wire 1 [? outputLine $end
$var wire 2 p? selectLines [1:0] $end
$var wire 2 q? w [1:0] $end
$scope module M0 $end
$var wire 2 r? inputLines [1:0] $end
$var wire 1 s? outputLine $end
$var wire 1 t? selectLine $end
$var wire 1 u? w1 $end
$var wire 1 v? w2 $end
$var wire 1 w? w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 x? inputLines [1:0] $end
$var wire 1 y? outputLine $end
$var wire 1 z? selectLine $end
$var wire 1 {? w1 $end
$var wire 1 |? w2 $end
$var wire 1 }? w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 ~? inputLines [1:0] $end
$var wire 1 [? outputLine $end
$var wire 1 !@ selectLine $end
$var wire 1 "@ w1 $end
$var wire 1 #@ w2 $end
$var wire 1 $@ w3 $end
$upscope $end
$upscope $end
$upscope $end
$scope module A63 $end
$var wire 1 %@ Ainvert $end
$var wire 1 &@ Binvert $end
$var wire 1 '@ CarryIn $end
$var wire 1 (@ CarryOut $end
$var wire 1 )@ Less $end
$var wire 2 *@ Operation [1:0] $end
$var wire 1 " Overflow $end
$var wire 1 +@ Result $end
$var wire 1 3 Set $end
$var wire 1 ,@ a $end
$var wire 1 -@ b $end
$var wire 2 .@ mux0inputs [1:0] $end
$var wire 2 /@ mux1inputs [1:0] $end
$var wire 4 0@ mux2inputs [3:0] $end
$var wire 1 1@ w1 $end
$var wire 1 2@ w2 $end
$scope module J0 $end
$var wire 2 3@ inputLines [1:0] $end
$var wire 1 1@ outputLine $end
$var wire 1 %@ selectLine $end
$var wire 1 4@ w1 $end
$var wire 1 5@ w2 $end
$var wire 1 6@ w3 $end
$upscope $end
$scope module J1 $end
$var wire 2 7@ inputLines [1:0] $end
$var wire 1 2@ outputLine $end
$var wire 1 &@ selectLine $end
$var wire 1 8@ w1 $end
$var wire 1 9@ w2 $end
$var wire 1 :@ w3 $end
$upscope $end
$scope module fa0 $end
$var wire 1 1@ a $end
$var wire 1 2@ b $end
$var wire 1 '@ cin $end
$var wire 1 (@ cout $end
$var wire 1 ;@ sum $end
$var wire 1 <@ w1 $end
$var wire 1 =@ w2 $end
$var wire 1 >@ w3 $end
$upscope $end
$scope module J5 $end
$var wire 4 ?@ inputLines [3:0] $end
$var wire 1 +@ outputLine $end
$var wire 2 @@ selectLines [1:0] $end
$var wire 2 A@ w [1:0] $end
$scope module M0 $end
$var wire 2 B@ inputLines [1:0] $end
$var wire 1 C@ outputLine $end
$var wire 1 D@ selectLine $end
$var wire 1 E@ w1 $end
$var wire 1 F@ w2 $end
$var wire 1 G@ w3 $end
$upscope $end
$scope module M1 $end
$var wire 2 H@ inputLines [1:0] $end
$var wire 1 I@ outputLine $end
$var wire 1 J@ selectLine $end
$var wire 1 K@ w1 $end
$var wire 1 L@ w2 $end
$var wire 1 M@ w3 $end
$upscope $end
$scope module M2 $end
$var wire 2 N@ inputLines [1:0] $end
$var wire 1 +@ outputLine $end
$var wire 1 O@ selectLine $end
$var wire 1 P@ w1 $end
$var wire 1 Q@ w2 $end
$var wire 1 R@ w3 $end
$upscope $end
$upscope $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
xR@
xQ@
xP@
xO@
bx N@
0M@
xL@
xK@
xJ@
xI@
b0x H@
xG@
xF@
xE@
xD@
xC@
bx B@
bx A@
bx @@
b0xxx ?@
x>@
x=@
x<@
x;@
x:@
x9@
x8@
bx 7@
x6@
x5@
x4@
bx 3@
x2@
x1@
b0xxx 0@
bx /@
bx .@
x-@
x,@
x+@
bx *@
0)@
x(@
x'@
x&@
x%@
x$@
x#@
x"@
x!@
bx ~?
0}?
x|?
x{?
xz?
xy?
b0x x?
xw?
xv?
xu?
xt?
xs?
bx r?
bx q?
bx p?
b0xxx o?
xn?
xm?
xl?
xk?
xj?
xi?
xh?
bx g?
xf?
xe?
xd?
bx c?
xb?
xa?
b0xxx `?
bx _?
bx ^?
x]?
x\?
x[?
bx Z?
0Y?
xX?
xW?
xV?
xU?
xT?
xS?
xR?
xQ?
bx P?
0O?
xN?
xM?
xL?
xK?
b0x J?
xI?
xH?
xG?
xF?
xE?
bx D?
bx C?
bx B?
b0xxx A?
x@?
x??
x>?
x=?
x<?
x;?
x:?
bx 9?
x8?
x7?
x6?
bx 5?
x4?
x3?
b0xxx 2?
bx 1?
bx 0?
x/?
x.?
x-?
bx ,?
0+?
x*?
x)?
x(?
x'?
x&?
x%?
x$?
x#?
bx "?
0!?
x~>
x}>
x|>
x{>
b0x z>
xy>
xx>
xw>
xv>
xu>
bx t>
bx s>
bx r>
b0xxx q>
xp>
xo>
xn>
xm>
xl>
xk>
xj>
bx i>
xh>
xg>
xf>
bx e>
xd>
xc>
b0xxx b>
bx a>
bx `>
x_>
x^>
x]>
bx \>
0[>
xZ>
xY>
xX>
xW>
xV>
xU>
xT>
xS>
bx R>
0Q>
xP>
xO>
xN>
xM>
b0x L>
xK>
xJ>
xI>
xH>
xG>
bx F>
bx E>
bx D>
b0xxx C>
xB>
xA>
x@>
x?>
x>>
x=>
x<>
bx ;>
x:>
x9>
x8>
bx 7>
x6>
x5>
b0xxx 4>
bx 3>
bx 2>
x1>
x0>
x/>
bx .>
0->
x,>
x+>
x*>
x)>
x(>
x'>
x&>
x%>
bx $>
0#>
x">
x!>
x~=
x}=
b0x |=
x{=
xz=
xy=
xx=
xw=
bx v=
bx u=
bx t=
b0xxx s=
xr=
xq=
xp=
xo=
xn=
xm=
xl=
bx k=
xj=
xi=
xh=
bx g=
xf=
xe=
b0xxx d=
bx c=
bx b=
xa=
x`=
x_=
bx ^=
0]=
x\=
x[=
xZ=
xY=
xX=
xW=
xV=
xU=
bx T=
0S=
xR=
xQ=
xP=
xO=
b0x N=
xM=
xL=
xK=
xJ=
xI=
bx H=
bx G=
bx F=
b0xxx E=
xD=
xC=
xB=
xA=
x@=
x?=
x>=
bx ==
x<=
x;=
x:=
bx 9=
x8=
x7=
b0xxx 6=
bx 5=
bx 4=
x3=
x2=
x1=
bx 0=
0/=
x.=
x-=
x,=
x+=
x*=
x)=
x(=
x'=
bx &=
0%=
x$=
x#=
x"=
x!=
b0x ~<
x}<
x|<
x{<
xz<
xy<
bx x<
bx w<
bx v<
b0xxx u<
xt<
xs<
xr<
xq<
xp<
xo<
xn<
bx m<
xl<
xk<
xj<
bx i<
xh<
xg<
b0xxx f<
bx e<
bx d<
xc<
xb<
xa<
bx `<
0_<
x^<
x]<
x\<
x[<
xZ<
xY<
xX<
xW<
bx V<
0U<
xT<
xS<
xR<
xQ<
b0x P<
xO<
xN<
xM<
xL<
xK<
bx J<
bx I<
bx H<
b0xxx G<
xF<
xE<
xD<
xC<
xB<
xA<
x@<
bx ?<
x><
x=<
x<<
bx ;<
x:<
x9<
b0xxx 8<
bx 7<
bx 6<
x5<
x4<
x3<
bx 2<
01<
x0<
x/<
x.<
x-<
x,<
x+<
x*<
x)<
bx (<
0'<
x&<
x%<
x$<
x#<
b0x "<
x!<
x~;
x};
x|;
x{;
bx z;
bx y;
bx x;
b0xxx w;
xv;
xu;
xt;
xs;
xr;
xq;
xp;
bx o;
xn;
xm;
xl;
bx k;
xj;
xi;
b0xxx h;
bx g;
bx f;
xe;
xd;
xc;
bx b;
0a;
x`;
x_;
x^;
x];
x\;
x[;
xZ;
xY;
bx X;
0W;
xV;
xU;
xT;
xS;
b0x R;
xQ;
xP;
xO;
xN;
xM;
bx L;
bx K;
bx J;
b0xxx I;
xH;
xG;
xF;
xE;
xD;
xC;
xB;
bx A;
x@;
x?;
x>;
bx =;
x<;
x;;
b0xxx :;
bx 9;
bx 8;
x7;
x6;
x5;
bx 4;
03;
x2;
x1;
x0;
x/;
x.;
x-;
x,;
x+;
bx *;
0);
x(;
x';
x&;
x%;
b0x $;
x#;
x";
x!;
x~:
x}:
bx |:
bx {:
bx z:
b0xxx y:
xx:
xw:
xv:
xu:
xt:
xs:
xr:
bx q:
xp:
xo:
xn:
bx m:
xl:
xk:
b0xxx j:
bx i:
bx h:
xg:
xf:
xe:
bx d:
0c:
xb:
xa:
x`:
x_:
x^:
x]:
x\:
x[:
bx Z:
0Y:
xX:
xW:
xV:
xU:
b0x T:
xS:
xR:
xQ:
xP:
xO:
bx N:
bx M:
bx L:
b0xxx K:
xJ:
xI:
xH:
xG:
xF:
xE:
xD:
bx C:
xB:
xA:
x@:
bx ?:
x>:
x=:
b0xxx <:
bx ;:
bx ::
x9:
x8:
x7:
bx 6:
05:
x4:
x3:
x2:
x1:
x0:
x/:
x.:
x-:
bx ,:
0+:
x*:
x):
x(:
x':
b0x &:
x%:
x$:
x#:
x":
x!:
bx ~9
bx }9
bx |9
b0xxx {9
xz9
xy9
xx9
xw9
xv9
xu9
xt9
bx s9
xr9
xq9
xp9
bx o9
xn9
xm9
b0xxx l9
bx k9
bx j9
xi9
xh9
xg9
bx f9
0e9
xd9
xc9
xb9
xa9
x`9
x_9
x^9
x]9
bx \9
0[9
xZ9
xY9
xX9
xW9
b0x V9
xU9
xT9
xS9
xR9
xQ9
bx P9
bx O9
bx N9
b0xxx M9
xL9
xK9
xJ9
xI9
xH9
xG9
xF9
bx E9
xD9
xC9
xB9
bx A9
x@9
x?9
b0xxx >9
bx =9
bx <9
x;9
x:9
x99
bx 89
079
x69
x59
x49
x39
x29
x19
x09
x/9
bx .9
0-9
x,9
x+9
x*9
x)9
b0x (9
x'9
x&9
x%9
x$9
x#9
bx "9
bx !9
bx ~8
b0xxx }8
x|8
x{8
xz8
xy8
xx8
xw8
xv8
bx u8
xt8
xs8
xr8
bx q8
xp8
xo8
b0xxx n8
bx m8
bx l8
xk8
xj8
xi8
bx h8
0g8
xf8
xe8
xd8
xc8
xb8
xa8
x`8
x_8
bx ^8
0]8
x\8
x[8
xZ8
xY8
b0x X8
xW8
xV8
xU8
xT8
xS8
bx R8
bx Q8
bx P8
b0xxx O8
xN8
xM8
xL8
xK8
xJ8
xI8
xH8
bx G8
xF8
xE8
xD8
bx C8
xB8
xA8
b0xxx @8
bx ?8
bx >8
x=8
x<8
x;8
bx :8
098
x88
x78
x68
x58
x48
x38
x28
x18
bx 08
0/8
x.8
x-8
x,8
x+8
b0x *8
x)8
x(8
x'8
x&8
x%8
bx $8
bx #8
bx "8
b0xxx !8
x~7
x}7
x|7
x{7
xz7
xy7
xx7
bx w7
xv7
xu7
xt7
bx s7
xr7
xq7
b0xxx p7
bx o7
bx n7
xm7
xl7
xk7
bx j7
0i7
xh7
xg7
xf7
xe7
xd7
xc7
xb7
xa7
bx `7
0_7
x^7
x]7
x\7
x[7
b0x Z7
xY7
xX7
xW7
xV7
xU7
bx T7
bx S7
bx R7
b0xxx Q7
xP7
xO7
xN7
xM7
xL7
xK7
xJ7
bx I7
xH7
xG7
xF7
bx E7
xD7
xC7
b0xxx B7
bx A7
bx @7
x?7
x>7
x=7
bx <7
0;7
x:7
x97
x87
x77
x67
x57
x47
x37
bx 27
017
x07
x/7
x.7
x-7
b0x ,7
x+7
x*7
x)7
x(7
x'7
bx &7
bx %7
bx $7
b0xxx #7
x"7
x!7
x~6
x}6
x|6
x{6
xz6
bx y6
xx6
xw6
xv6
bx u6
xt6
xs6
b0xxx r6
bx q6
bx p6
xo6
xn6
xm6
bx l6
0k6
xj6
xi6
xh6
xg6
xf6
xe6
xd6
xc6
bx b6
0a6
x`6
x_6
x^6
x]6
b0x \6
x[6
xZ6
xY6
xX6
xW6
bx V6
bx U6
bx T6
b0xxx S6
xR6
xQ6
xP6
xO6
xN6
xM6
xL6
bx K6
xJ6
xI6
xH6
bx G6
xF6
xE6
b0xxx D6
bx C6
bx B6
xA6
x@6
x?6
bx >6
0=6
x<6
x;6
x:6
x96
x86
x76
x66
x56
bx 46
036
x26
x16
x06
x/6
b0x .6
x-6
x,6
x+6
x*6
x)6
bx (6
bx '6
bx &6
b0xxx %6
x$6
x#6
x"6
x!6
x~5
x}5
x|5
bx {5
xz5
xy5
xx5
bx w5
xv5
xu5
b0xxx t5
bx s5
bx r5
xq5
xp5
xo5
bx n5
0m5
xl5
xk5
xj5
xi5
xh5
xg5
xf5
xe5
bx d5
0c5
xb5
xa5
x`5
x_5
b0x ^5
x]5
x\5
x[5
xZ5
xY5
bx X5
bx W5
bx V5
b0xxx U5
xT5
xS5
xR5
xQ5
xP5
xO5
xN5
bx M5
xL5
xK5
xJ5
bx I5
xH5
xG5
b0xxx F5
bx E5
bx D5
xC5
xB5
xA5
bx @5
0?5
x>5
x=5
x<5
x;5
x:5
x95
x85
x75
bx 65
055
x45
x35
x25
x15
b0x 05
x/5
x.5
x-5
x,5
x+5
bx *5
bx )5
bx (5
b0xxx '5
x&5
x%5
x$5
x#5
x"5
x!5
x~4
bx }4
x|4
x{4
xz4
bx y4
xx4
xw4
b0xxx v4
bx u4
bx t4
xs4
xr4
xq4
bx p4
0o4
xn4
xm4
xl4
xk4
xj4
xi4
xh4
xg4
bx f4
0e4
xd4
xc4
xb4
xa4
b0x `4
x_4
x^4
x]4
x\4
x[4
bx Z4
bx Y4
bx X4
b0xxx W4
xV4
xU4
xT4
xS4
xR4
xQ4
xP4
bx O4
xN4
xM4
xL4
bx K4
xJ4
xI4
b0xxx H4
bx G4
bx F4
xE4
xD4
xC4
bx B4
0A4
x@4
x?4
x>4
x=4
x<4
x;4
x:4
x94
bx 84
074
x64
x54
x44
x34
b0x 24
x14
x04
x/4
x.4
x-4
bx ,4
bx +4
bx *4
b0xxx )4
x(4
x'4
x&4
x%4
x$4
x#4
x"4
bx !4
x~3
x}3
x|3
bx {3
xz3
xy3
b0xxx x3
bx w3
bx v3
xu3
xt3
xs3
bx r3
0q3
xp3
xo3
xn3
xm3
xl3
xk3
xj3
xi3
bx h3
0g3
xf3
xe3
xd3
xc3
b0x b3
xa3
x`3
x_3
x^3
x]3
bx \3
bx [3
bx Z3
b0xxx Y3
xX3
xW3
xV3
xU3
xT3
xS3
xR3
bx Q3
xP3
xO3
xN3
bx M3
xL3
xK3
b0xxx J3
bx I3
bx H3
xG3
xF3
xE3
bx D3
0C3
xB3
xA3
x@3
x?3
x>3
x=3
x<3
x;3
bx :3
093
x83
x73
x63
x53
b0x 43
x33
x23
x13
x03
x/3
bx .3
bx -3
bx ,3
b0xxx +3
x*3
x)3
x(3
x'3
x&3
x%3
x$3
bx #3
x"3
x!3
x~2
bx }2
x|2
x{2
b0xxx z2
bx y2
bx x2
xw2
xv2
xu2
bx t2
0s2
xr2
xq2
xp2
xo2
xn2
xm2
xl2
xk2
bx j2
0i2
xh2
xg2
xf2
xe2
b0x d2
xc2
xb2
xa2
x`2
x_2
bx ^2
bx ]2
bx \2
b0xxx [2
xZ2
xY2
xX2
xW2
xV2
xU2
xT2
bx S2
xR2
xQ2
xP2
bx O2
xN2
xM2
b0xxx L2
bx K2
bx J2
xI2
xH2
xG2
bx F2
0E2
xD2
xC2
xB2
xA2
x@2
x?2
x>2
x=2
bx <2
0;2
x:2
x92
x82
x72
b0x 62
x52
x42
x32
x22
x12
bx 02
bx /2
bx .2
b0xxx -2
x,2
x+2
x*2
x)2
x(2
x'2
x&2
bx %2
x$2
x#2
x"2
bx !2
x~1
x}1
b0xxx |1
bx {1
bx z1
xy1
xx1
xw1
bx v1
0u1
xt1
xs1
xr1
xq1
xp1
xo1
xn1
xm1
bx l1
0k1
xj1
xi1
xh1
xg1
b0x f1
xe1
xd1
xc1
xb1
xa1
bx `1
bx _1
bx ^1
b0xxx ]1
x\1
x[1
xZ1
xY1
xX1
xW1
xV1
bx U1
xT1
xS1
xR1
bx Q1
xP1
xO1
b0xxx N1
bx M1
bx L1
xK1
xJ1
xI1
bx H1
0G1
xF1
xE1
xD1
xC1
xB1
xA1
x@1
x?1
bx >1
0=1
x<1
x;1
x:1
x91
b0x 81
x71
x61
x51
x41
x31
bx 21
bx 11
bx 01
b0xxx /1
x.1
x-1
x,1
x+1
x*1
x)1
x(1
bx '1
x&1
x%1
x$1
bx #1
x"1
x!1
b0xxx ~0
bx }0
bx |0
x{0
xz0
xy0
bx x0
0w0
xv0
xu0
xt0
xs0
xr0
xq0
xp0
xo0
bx n0
0m0
xl0
xk0
xj0
xi0
b0x h0
xg0
xf0
xe0
xd0
xc0
bx b0
bx a0
bx `0
b0xxx _0
x^0
x]0
x\0
x[0
xZ0
xY0
xX0
bx W0
xV0
xU0
xT0
bx S0
xR0
xQ0
b0xxx P0
bx O0
bx N0
xM0
xL0
xK0
bx J0
0I0
xH0
xG0
xF0
xE0
xD0
xC0
xB0
xA0
bx @0
0?0
x>0
x=0
x<0
x;0
b0x :0
x90
x80
x70
x60
x50
bx 40
bx 30
bx 20
b0xxx 10
x00
x/0
x.0
x-0
x,0
x+0
x*0
bx )0
x(0
x'0
x&0
bx %0
x$0
x#0
b0xxx "0
bx !0
bx ~/
x}/
x|/
x{/
bx z/
0y/
xx/
xw/
xv/
xu/
xt/
xs/
xr/
xq/
bx p/
0o/
xn/
xm/
xl/
xk/
b0x j/
xi/
xh/
xg/
xf/
xe/
bx d/
bx c/
bx b/
b0xxx a/
x`/
x_/
x^/
x]/
x\/
x[/
xZ/
bx Y/
xX/
xW/
xV/
bx U/
xT/
xS/
b0xxx R/
bx Q/
bx P/
xO/
xN/
xM/
bx L/
0K/
xJ/
xI/
xH/
xG/
xF/
xE/
xD/
xC/
bx B/
0A/
x@/
x?/
x>/
x=/
b0x </
x;/
x:/
x9/
x8/
x7/
bx 6/
bx 5/
bx 4/
b0xxx 3/
x2/
x1/
x0/
x//
x./
x-/
x,/
bx +/
x*/
x)/
x(/
bx '/
x&/
x%/
b0xxx $/
bx #/
bx "/
x!/
x~.
x}.
bx |.
0{.
xz.
xy.
xx.
xw.
xv.
xu.
xt.
xs.
bx r.
0q.
xp.
xo.
xn.
xm.
b0x l.
xk.
xj.
xi.
xh.
xg.
bx f.
bx e.
bx d.
b0xxx c.
xb.
xa.
x`.
x_.
x^.
x].
x\.
bx [.
xZ.
xY.
xX.
bx W.
xV.
xU.
b0xxx T.
bx S.
bx R.
xQ.
xP.
xO.
bx N.
0M.
xL.
xK.
xJ.
xI.
xH.
xG.
xF.
xE.
bx D.
0C.
xB.
xA.
x@.
x?.
b0x >.
x=.
x<.
x;.
x:.
x9.
bx 8.
bx 7.
bx 6.
b0xxx 5.
x4.
x3.
x2.
x1.
x0.
x/.
x..
bx -.
x,.
x+.
x*.
bx ).
x(.
x'.
b0xxx &.
bx %.
bx $.
x#.
x".
x!.
bx ~-
0}-
x|-
x{-
xz-
xy-
xx-
xw-
xv-
xu-
bx t-
0s-
xr-
xq-
xp-
xo-
b0x n-
xm-
xl-
xk-
xj-
xi-
bx h-
bx g-
bx f-
b0xxx e-
xd-
xc-
xb-
xa-
x`-
x_-
x^-
bx ]-
x\-
x[-
xZ-
bx Y-
xX-
xW-
b0xxx V-
bx U-
bx T-
xS-
xR-
xQ-
bx P-
0O-
xN-
xM-
xL-
xK-
xJ-
xI-
xH-
xG-
bx F-
0E-
xD-
xC-
xB-
xA-
b0x @-
x?-
x>-
x=-
x<-
x;-
bx :-
bx 9-
bx 8-
b0xxx 7-
x6-
x5-
x4-
x3-
x2-
x1-
x0-
bx /-
x.-
x--
x,-
bx +-
x*-
x)-
b0xxx (-
bx '-
bx &-
x%-
x$-
x#-
bx "-
0!-
x~,
x},
x|,
x{,
xz,
xy,
xx,
xw,
bx v,
0u,
xt,
xs,
xr,
xq,
b0x p,
xo,
xn,
xm,
xl,
xk,
bx j,
bx i,
bx h,
b0xxx g,
xf,
xe,
xd,
xc,
xb,
xa,
x`,
bx _,
x^,
x],
x\,
bx [,
xZ,
xY,
b0xxx X,
bx W,
bx V,
xU,
xT,
xS,
bx R,
0Q,
xP,
xO,
xN,
xM,
xL,
xK,
xJ,
xI,
bx H,
0G,
xF,
xE,
xD,
xC,
b0x B,
xA,
x@,
x?,
x>,
x=,
bx <,
bx ;,
bx :,
b0xxx 9,
x8,
x7,
x6,
x5,
x4,
x3,
x2,
bx 1,
x0,
x/,
x.,
bx -,
x,,
x+,
b0xxx *,
bx ),
bx (,
x',
x&,
x%,
bx $,
0#,
x",
x!,
x~+
x}+
x|+
x{+
xz+
xy+
bx x+
0w+
xv+
xu+
xt+
xs+
b0x r+
xq+
xp+
xo+
xn+
xm+
bx l+
bx k+
bx j+
b0xxx i+
xh+
xg+
xf+
xe+
xd+
xc+
xb+
bx a+
x`+
x_+
x^+
bx ]+
x\+
x[+
b0xxx Z+
bx Y+
bx X+
xW+
xV+
xU+
bx T+
0S+
xR+
xQ+
xP+
xO+
xN+
xM+
xL+
xK+
bx J+
0I+
xH+
xG+
xF+
xE+
b0x D+
xC+
xB+
xA+
x@+
x?+
bx >+
bx =+
bx <+
b0xxx ;+
x:+
x9+
x8+
x7+
x6+
x5+
x4+
bx 3+
x2+
x1+
x0+
bx /+
x.+
x-+
b0xxx ,+
bx ++
bx *+
x)+
x(+
x'+
bx &+
0%+
x$+
x#+
x"+
x!+
x~*
x}*
x|*
x{*
bx z*
0y*
xx*
xw*
xv*
xu*
b0x t*
xs*
xr*
xq*
xp*
xo*
bx n*
bx m*
bx l*
b0xxx k*
xj*
xi*
xh*
xg*
xf*
xe*
xd*
bx c*
xb*
xa*
x`*
bx _*
x^*
x]*
b0xxx \*
bx [*
bx Z*
xY*
xX*
xW*
bx V*
0U*
xT*
xS*
xR*
xQ*
xP*
xO*
xN*
xM*
bx L*
0K*
xJ*
xI*
xH*
xG*
b0x F*
xE*
xD*
xC*
xB*
xA*
bx @*
bx ?*
bx >*
b0xxx =*
x<*
x;*
x:*
x9*
x8*
x7*
x6*
bx 5*
x4*
x3*
x2*
bx 1*
x0*
x/*
b0xxx .*
bx -*
bx ,*
x+*
x**
x)*
bx (*
0'*
x&*
x%*
x$*
x#*
x"*
x!*
x~)
x})
bx |)
0{)
xz)
xy)
xx)
xw)
b0x v)
xu)
xt)
xs)
xr)
xq)
bx p)
bx o)
bx n)
b0xxx m)
xl)
xk)
xj)
xi)
xh)
xg)
xf)
bx e)
xd)
xc)
xb)
bx a)
x`)
x_)
b0xxx ^)
bx ])
bx \)
x[)
xZ)
xY)
bx X)
0W)
xV)
xU)
xT)
xS)
xR)
xQ)
xP)
xO)
bx N)
0M)
xL)
xK)
xJ)
xI)
b0x H)
xG)
xF)
xE)
xD)
xC)
bx B)
bx A)
bx @)
b0xxx ?)
x>)
x=)
x<)
x;)
x:)
x9)
x8)
bx 7)
x6)
x5)
x4)
bx 3)
x2)
x1)
b0xxx 0)
bx /)
bx .)
x-)
x,)
x+)
bx *)
0))
x()
x')
x&)
x%)
x$)
x#)
x")
x!)
bx ~(
0}(
x|(
x{(
xz(
xy(
b0x x(
xw(
xv(
xu(
xt(
xs(
bx r(
bx q(
bx p(
b0xxx o(
xn(
xm(
xl(
xk(
xj(
xi(
xh(
bx g(
xf(
xe(
xd(
bx c(
xb(
xa(
b0xxx `(
bx _(
bx ^(
x](
x\(
x[(
bx Z(
0Y(
xX(
xW(
xV(
xU(
xT(
xS(
xR(
xQ(
bx P(
0O(
xN(
xM(
xL(
xK(
b0x J(
xI(
xH(
xG(
xF(
xE(
bx D(
bx C(
bx B(
b0xxx A(
x@(
x?(
x>(
x=(
x<(
x;(
x:(
bx 9(
x8(
x7(
x6(
bx 5(
x4(
x3(
b0xxx 2(
bx 1(
bx 0(
x/(
x.(
x-(
bx ,(
0+(
x*(
x)(
x((
x'(
x&(
x%(
x$(
x#(
bx "(
0!(
x~'
x}'
x|'
x{'
b0x z'
xy'
xx'
xw'
xv'
xu'
bx t'
bx s'
bx r'
b0xxx q'
xp'
xo'
xn'
xm'
xl'
xk'
xj'
bx i'
xh'
xg'
xf'
bx e'
xd'
xc'
b0xxx b'
bx a'
bx `'
x_'
x^'
x]'
bx \'
0['
xZ'
xY'
xX'
xW'
xV'
xU'
xT'
xS'
bx R'
0Q'
xP'
xO'
xN'
xM'
b0x L'
xK'
xJ'
xI'
xH'
xG'
bx F'
bx E'
bx D'
b0xxx C'
xB'
xA'
x@'
x?'
x>'
x='
x<'
bx ;'
x:'
x9'
x8'
bx 7'
x6'
x5'
b0xxx 4'
bx 3'
bx 2'
x1'
x0'
x/'
bx .'
0-'
x,'
x+'
x*'
x)'
x('
x''
x&'
x%'
bx $'
0#'
x"'
x!'
x~&
x}&
b0x |&
x{&
xz&
xy&
xx&
xw&
bx v&
bx u&
bx t&
b0xxx s&
xr&
xq&
xp&
xo&
xn&
xm&
xl&
bx k&
xj&
xi&
xh&
bx g&
xf&
xe&
b0xxx d&
bx c&
bx b&
xa&
x`&
x_&
bx ^&
0]&
x\&
x[&
xZ&
xY&
xX&
xW&
xV&
xU&
bx T&
0S&
xR&
xQ&
xP&
xO&
b0x N&
xM&
xL&
xK&
xJ&
xI&
bx H&
bx G&
bx F&
b0xxx E&
xD&
xC&
xB&
xA&
x@&
x?&
x>&
bx =&
x<&
x;&
x:&
bx 9&
x8&
x7&
b0xxx 6&
bx 5&
bx 4&
x3&
x2&
x1&
bx 0&
0/&
x.&
x-&
x,&
x+&
x*&
x)&
x(&
x'&
bx &&
0%&
x$&
x#&
x"&
x!&
b0x ~%
x}%
x|%
x{%
xz%
xy%
bx x%
bx w%
bx v%
b0xxx u%
xt%
xs%
xr%
xq%
xp%
xo%
xn%
bx m%
xl%
xk%
xj%
bx i%
xh%
xg%
b0xxx f%
bx e%
bx d%
xc%
xb%
xa%
bx `%
0_%
x^%
x]%
x\%
x[%
xZ%
xY%
xX%
xW%
bx V%
0U%
xT%
xS%
xR%
xQ%
b0x P%
xO%
xN%
xM%
xL%
xK%
bx J%
bx I%
bx H%
b0xxx G%
xF%
xE%
xD%
xC%
xB%
xA%
x@%
bx ?%
x>%
x=%
x<%
bx ;%
x:%
x9%
b0xxx 8%
bx 7%
bx 6%
x5%
x4%
x3%
bx 2%
01%
x0%
x/%
x.%
x-%
x,%
x+%
x*%
x)%
bx (%
0'%
x&%
x%%
x$%
x#%
b0x "%
x!%
x~$
x}$
x|$
x{$
bx z$
bx y$
bx x$
b0xxx w$
xv$
xu$
xt$
xs$
xr$
xq$
xp$
bx o$
xn$
xm$
xl$
bx k$
xj$
xi$
b0xxx h$
bx g$
bx f$
xe$
xd$
xc$
bx b$
0a$
x`$
x_$
x^$
x]$
x\$
x[$
xZ$
xY$
bx X$
0W$
xV$
xU$
xT$
xS$
b0x R$
xQ$
xP$
xO$
xN$
xM$
bx L$
bx K$
bx J$
b0xxx I$
xH$
xG$
xF$
xE$
xD$
xC$
xB$
bx A$
x@$
x?$
x>$
bx =$
x<$
x;$
b0xxx :$
bx 9$
bx 8$
x7$
x6$
x5$
bx 4$
03$
x2$
x1$
x0$
x/$
x.$
x-$
x,$
x+$
bx *$
0)$
x($
x'$
x&$
x%$
b0x $$
x#$
x"$
x!$
x~#
x}#
bx |#
bx {#
bx z#
b0xxx y#
xx#
xw#
xv#
xu#
xt#
xs#
xr#
bx q#
xp#
xo#
xn#
bx m#
xl#
xk#
b0xxx j#
bx i#
bx h#
xg#
xf#
xe#
bx d#
0c#
xb#
xa#
x`#
x_#
x^#
x]#
x\#
x[#
bx Z#
0Y#
xX#
xW#
xV#
xU#
b0x T#
xS#
xR#
xQ#
xP#
xO#
bx N#
bx M#
bx L#
b0xxx K#
xJ#
xI#
xH#
xG#
xF#
xE#
xD#
bx C#
xB#
xA#
x@#
bx ?#
x>#
x=#
b0xxx <#
bx ;#
bx :#
x9#
x8#
x7#
bx 6#
05#
x4#
x3#
x2#
x1#
x0#
x/#
x.#
x-#
bx ,#
0+#
x*#
x)#
x(#
x'#
b0x &#
x%#
x$#
x##
x"#
x!#
bx ~"
bx }"
bx |"
b0xxx {"
xz"
xy"
xx"
xw"
xv"
xu"
xt"
bx s"
xr"
xq"
xp"
bx o"
xn"
xm"
b0xxx l"
bx k"
bx j"
xi"
xh"
xg"
bx f"
0e"
xd"
xc"
xb"
xa"
x`"
x_"
x^"
x]"
bx \"
0["
xZ"
xY"
xX"
xW"
b0x V"
xU"
xT"
xS"
xR"
xQ"
bx P"
bx O"
bx N"
b0xxx M"
xL"
xK"
xJ"
xI"
xH"
xG"
xF"
bx E"
xD"
xC"
xB"
bx A"
x@"
x?"
b0xxx >"
bx ="
bx <"
x;"
x:"
x9"
bx 8"
07"
x6"
x5"
x4"
x3"
x2"
x1"
x0"
x/"
bx ."
0-"
x,"
x+"
x*"
x)"
b0x ("
x'"
x&"
x%"
x$"
x#"
bx ""
bx !"
bx ~
b0xxx }
x|
x{
xz
xy
xx
xw
xv
bx u
xt
xs
xr
bx q
xp
xo
b0xxx n
bx m
bx l
xk
xj
xi
bx h
0g
xf
xe
xd
xc
xb
xa
x`
x_
bx ^
x]
x\
x[
xZ
xY
bx X
xW
xV
xU
xT
xS
bx R
bx Q
bx P
bx O
xN
xM
xL
xK
xJ
xI
xH
bx G
xF
xE
xD
bx C
xB
xA
bx @
bx ?
bx >
x=
x<
x;
bx :
x9
x8
x7
x6
bx 5
bx 4
x3
bx 2
bx 1
bx 0
bx /
bx .
bx -
bx ,
bx +
bx *
bx )
bx (
bx '
bx &
bx %
x$
bx #
x"
bx !
$end
#5
0$
0%$
0!&
0($
0$&
1)"
1;
0W"
0'#
1U#
b0 $$
0S$
0#%
1Q%
b0 ~%
0O&
0}&
0M'
0{'
0K(
0y(
0I)
0w)
0G*
0u*
0E+
0s+
0C,
0q,
0A-
0o-
0?.
0m.
0Y8
0=/
0}=
0k/
0;0
0i0
091
0g1
072
0e2
053
0c3
034
0a4
015
0_5
0/6
0]6
0-7
0[7
0+8
0)9
0W9
0':
0U:
0%;
0S;
0#<
0Q<
0!=
0O=
0M>
0{>
0K?
0y?
0I@
03%
1,"
1a
0Z"
0i
0*#
09"
1X#
0u#
0g"
07#
0V$
0e#
0&%
05$
1T%
0q%
0c$
0R&
0a%
0"'
01&
0P'
0_&
0~'
0/'
0N(
0]'
0|(
0-(
0L)
0[(
0z)
0+)
0J*
0Y)
0x*
0)*
0H+
0W*
0v+
0'+
0F,
0U+
0t,
0%,
0D-
0S,
0r-
0#-
0B.
0Q-
0p.
0\8
0!.
0@/
0">
0O.
0n/
0}.
0>0
0M/
0l0
0{/
0<1
0K0
0j1
0y0
0:2
0I1
0h2
0w1
083
0G2
0f3
0u2
064
0E3
0d4
0s3
045
0C4
0b5
0q4
026
0A5
0`6
0o5
007
0?6
0^7
0m6
0.8
0=7
0k7
0,9
0;8
0Z9
0i8
0*:
099
0X:
0g9
0(;
07:
0V;
0e:
0&<
05;
0T<
0c;
0$=
03<
0R=
0a<
01=
0P>
0_=
0~>
0/>
0N?
0]>
0|?
0-?
0L@
0[?
0+@
b1 #
b1 2
0Y%
0Y
01"
0_"
0a#
0/#
0]#
0-$
0[$
0]%
0+%
0)&
0W&
0''
0U'
0%(
0S(
0#)
0Q)
0!*
0O*
0}*
0M+
0{+
0K,
0y,
0I-
0w-
0G.
0u.
0E/
0s/
0C0
0q0
0A1
0o1
0?2
0m2
0=3
0k3
0;4
0i4
095
0g5
076
0e6
057
0c7
038
0a8
019
0_9
0/:
0]:
0-;
0[;
0+<
0Y<
0)=
0W=
0'>
0U>
0%?
0S?
0#@
0Q@
0\
b1 ("
1S
b1 Q
b1 ^
b0 V"
b0 &#
b1 T#
04#
b0 R$
b0 "%
b1 P%
00%
b0 N&
b0 |&
b0 L'
b0 z'
b0 J(
b0 x(
b0 H)
b0 v)
b0 F*
b0 t*
b0 D+
b0 r+
b0 B,
b0 p,
b0 @-
b0 n-
b0 >.
b0 l.
b0 X8
b0 </
b0 |=
b0 j/
b0 :0
b0 h0
b0 81
b0 f1
b0 62
b0 d2
b0 43
b0 b3
b0 24
b0 `4
b0 05
b0 ^5
b0 .6
b0 \6
b0 ,7
b0 Z7
b0 *8
b0 (9
b0 V9
b0 &:
b0 T:
b0 $;
b0 R;
b0 "<
b0 P<
b0 ~<
b0 N=
b0 L>
b0 z>
b0 J?
b0 x?
03
b0 H@
0K%
b10 I%
b10 V%
1y
1V
0I"
0#"
b10 !"
b10 ."
0w"
0Q"
b0 O"
b0 \"
1G#
0J#
0!#
b0 }"
b0 ,#
0O#
b10 M#
b10 Z#
0E$
0}#
b0 {#
b0 *$
0s$
0M$
b0 K$
b0 X$
1C%
0F%
0{$
b0 y$
b0 (%
0A&
0y%
b0 w%
b0 &&
0o&
0I&
b0 G&
b0 T&
0?'
0w&
b0 u&
b0 $'
0m'
0G'
b0 E'
b0 R'
0=(
0u'
b0 s'
b0 "(
0k(
0E(
b0 C(
b0 P(
0;)
0s(
b0 q(
b0 ~(
0i)
0C)
b0 A)
b0 N)
09*
0q)
b0 o)
b0 |)
0g*
0A*
b0 ?*
b0 L*
07+
0o*
b0 m*
b0 z*
0e+
0?+
b0 =+
b0 J+
05,
0m+
b0 k+
b0 x+
0c,
0=,
b0 ;,
b0 H,
03-
0k,
b0 i,
b0 v,
0a-
0;-
b0 9-
b0 F-
01.
0i-
b0 g-
b0 t-
0_.
0K8
09.
b0 7.
b0 D.
0//
0o=
0g.
b0 e.
b0 r.
0]/
07/
b0 5/
b0 B/
0-0
0e/
b0 c/
b0 p/
0[0
050
b0 30
b0 @0
0+1
0c0
b0 a0
b0 n0
0Y1
031
b0 11
b0 >1
0)2
0a1
b0 _1
b0 l1
0W2
012
b0 /2
b0 <2
0'3
0_2
b0 ]2
b0 j2
0U3
0/3
b0 -3
b0 :3
0%4
0]3
b0 [3
b0 h3
0S4
0-4
b0 +4
b0 84
0#5
0[4
b0 Y4
b0 f4
0Q5
0+5
b0 )5
b0 65
0!6
0Y5
b0 W5
b0 d5
0O6
0)6
b0 '6
b0 46
0}6
0W6
b0 U6
b0 b6
0M7
0'7
b0 %7
b0 27
0{7
0U7
b0 S7
b0 `7
0%8
b0 #8
b0 08
0y8
0S8
b0 Q8
b0 ^8
0I9
0#9
b0 !9
b0 .9
0w9
0Q9
b0 O9
b0 \9
0G:
0!:
b0 }9
b0 ,:
0u:
0O:
b0 M:
b0 Z:
0E;
0}:
b0 {:
b0 *;
0s;
0M;
b0 K;
b0 X;
0C<
0{;
b0 y;
b0 (<
0q<
0K<
b0 I<
b0 V<
0A=
0y<
b0 w<
b0 &=
0I=
b0 G=
b0 T=
0?>
0w=
b0 u=
b0 $>
0m>
0G>
b0 E>
b0 R>
0=?
0u>
b0 s>
b0 "?
0k?
0E?
b0 C?
b0 P?
0"
0;@
0s?
b0 q?
b0 ~?
0C@
b0 A@
b0 N@
0N%
b0 X
1e
05"
0&"
0c"
0T"
03#
0$#
0R#
01$
0"$
0_$
0P$
0/%
0~$
0-&
0|%
0[&
0L&
0+'
0z&
0Y'
0J'
0)(
0x'
0W(
0H(
0')
0v(
0U)
0F)
0%*
0t)
0S*
0D*
0#+
0r*
0Q+
0B+
0!,
0p+
0O,
0@,
0},
0n,
0M-
0>-
0{-
0l-
0K.
078
0<.
0y.
0[=
0j.
0I/
0:/
0w/
0h/
0G0
080
0u0
0f0
0E1
061
0s1
0d1
0C2
042
0q2
0b2
0A3
023
0o3
0`3
0?4
004
0m4
0^4
0=5
0.5
0k5
0\5
0;6
0,6
0i6
0Z6
097
0*7
0g7
0X7
0(8
0e8
0V8
059
0&9
0c9
0T9
03:
0$:
0a:
0R:
01;
0";
0_;
0P;
0/<
0~;
0]<
0N<
0-=
0|<
0L=
0+>
0z=
0Y>
0J>
0)?
0x>
0W?
0H?
0'@
0v?
0F@
0K
19
b11 R
0f
06"
0d"
0b#
02$
0`$
0^%
0.&
0\&
0,'
0Z'
0*(
0X(
0()
0V)
0&*
0T*
0$+
0R+
0",
0P,
0~,
0N-
0|-
0L.
0z.
0J/
0x/
0H0
0v0
0F1
0t1
0D2
0r2
0B3
0p3
0@4
0n4
0>5
0l5
0<6
0j6
0:7
0h7
088
0f8
069
0d9
04:
0b:
02;
0`;
00<
0^<
0.=
0\=
0,>
0Z>
0*?
0X?
0(@
b1 1
1H#
b10 J%
0L
1M
b11 @
b11 O
0|
b0 ""
0L"
b0 P"
0z"
b0 ~"
b10 N#
0x#
b0 |#
0H$
b0 L$
0v$
b0 z$
0t%
b0 x%
0D&
b0 H&
0r&
b0 v&
0B'
b0 F'
0p'
b0 t'
0@(
b0 D(
0n(
b0 r(
0>)
b0 B)
0l)
b0 p)
0<*
b0 @*
0j*
b0 n*
0:+
b0 >+
0h+
b0 l+
08,
b0 <,
0f,
b0 j,
06-
b0 :-
0d-
b0 h-
04.
b0 8.
0b.
b0 f.
02/
b0 6/
0`/
b0 d/
000
b0 40
0^0
b0 b0
0.1
b0 21
0\1
b0 `1
0,2
b0 02
0Z2
b0 ^2
0*3
b0 .3
0X3
b0 \3
0(4
b0 ,4
0V4
b0 Z4
0&5
b0 *5
0T5
b0 X5
0$6
b0 (6
0R6
b0 V6
0"7
b0 &7
0P7
b0 T7
0~7
b0 $8
0N8
b0 R8
0|8
b0 "9
0L9
b0 P9
0z9
b0 ~9
0J:
b0 N:
0x:
b0 |:
0H;
b0 L;
0v;
b0 z;
0F<
b0 J<
0t<
b0 x<
0D=
b0 H=
0r=
b0 v=
0B>
b0 F>
0p>
b0 t>
0@?
b0 D?
0n?
b0 r?
0>@
b0 B@
1B
1>#
1D%
0E%
b110 8%
b110 G%
1A
0z
0{
b100 n
b100 }
0J"
0K"
b0 >"
b0 M"
0x"
0y"
b0 l"
b0 {"
0I#
b110 <#
b110 K#
0v#
0w#
b0 j#
b0 y#
0F$
0G$
b0 :$
b0 I$
0t$
0u$
b0 h$
b0 w$
19%
0r%
0s%
b0 f%
b0 u%
0B&
0C&
b0 6&
b0 E&
0p&
0q&
b0 d&
b0 s&
0@'
0A'
b0 4'
b0 C'
0n'
0o'
b0 b'
b0 q'
0>(
0?(
b0 2(
b0 A(
0l(
0m(
b0 `(
b0 o(
0<)
0=)
b0 0)
b0 ?)
0j)
0k)
b0 ^)
b0 m)
0:*
0;*
b0 .*
b0 =*
0h*
0i*
b0 \*
b0 k*
08+
09+
b0 ,+
b0 ;+
0f+
0g+
b0 Z+
b0 i+
06,
07,
b0 *,
b0 9,
0d,
0e,
b0 X,
b0 g,
04-
05-
b0 (-
b0 7-
0b-
0c-
b0 V-
b0 e-
02.
03.
b0 &.
b0 5.
0`.
0a.
b0 T.
b0 c.
00/
01/
b0 $/
b0 3/
0^/
0_/
b0 R/
b0 a/
0.0
0/0
b0 "0
b0 10
0\0
0]0
b0 P0
b0 _0
0,1
0-1
b0 ~0
b0 /1
0Z1
0[1
b0 N1
b0 ]1
0*2
0+2
b0 |1
b0 -2
0X2
0Y2
b0 L2
b0 [2
0(3
0)3
b0 z2
b0 +3
0V3
0W3
b0 J3
b0 Y3
0&4
0'4
b0 x3
b0 )4
0T4
0U4
b0 H4
b0 W4
0$5
0%5
b0 v4
b0 '5
0R5
0S5
b0 F5
b0 U5
0"6
0#6
b0 t5
b0 %6
0P6
0Q6
b0 D6
b0 S6
0~6
0!7
b0 r6
b0 #7
0N7
0O7
b0 B7
b0 Q7
0|7
0}7
b0 p7
b0 !8
0L8
0M8
b0 @8
b0 O8
0z8
0{8
b0 n8
b0 }8
0J9
0K9
b0 >9
b0 M9
0x9
0y9
b0 l9
b0 {9
0H:
0I:
b0 <:
b0 K:
0v:
0w:
b0 j:
b0 y:
0F;
0G;
b0 :;
b0 I;
0t;
0u;
b0 h;
b0 w;
0D<
0E<
b0 8<
b0 G<
0r<
0s<
b0 f<
b0 u<
0B=
0C=
b0 6=
b0 E=
0p=
0q=
b0 d=
b0 s=
0@>
0A>
b0 4>
b0 C>
0n>
0o>
b0 b>
b0 q>
0>?
0??
b0 2?
b0 A?
0l?
0m?
b0 `?
b0 o?
0<@
0=@
b0 0@
b0 ?@
1U
0W
1[
0]
1`
0b
1%"
0'"
1+"
10"
02"
1S"
0U"
1Y"
1^"
0`"
1##
0%#
1)#
1.#
00#
1Q#
0S#
1W#
1\#
0^#
1!$
0#$
1'$
1,$
0.$
1O$
0Q$
1U$
1Z$
0\$
1}$
0!%
1%%
1*%
0,%
1M%
0O%
1S%
1X%
0Z%
1{%
0}%
1#&
1(&
0*&
1K&
0M&
1Q&
1V&
0X&
1y&
0{&
1!'
1&'
0('
1I'
0K'
1O'
1T'
0V'
1w'
0y'
1}'
1$(
0&(
1G(
0I(
1M(
1R(
0T(
1u(
0w(
1{(
1")
0$)
1E)
0G)
1K)
1P)
0R)
1s)
0u)
1y)
1~)
0"*
1C*
0E*
1I*
1N*
0P*
1q*
0s*
1w*
1|*
0~*
1A+
0C+
1G+
1L+
0N+
1o+
0q+
1u+
1z+
0|+
1?,
0A,
1E,
1J,
0L,
1m,
0o,
1s,
1x,
0z,
1=-
0?-
1C-
1H-
0J-
1k-
0m-
1q-
1v-
0x-
1;.
0=.
1A.
1F.
0H.
1i.
0k.
1o.
1t.
0v.
19/
0;/
1?/
1D/
0F/
1g/
0i/
1m/
1r/
0t/
170
090
1=0
1B0
0D0
1e0
0g0
1k0
1p0
0r0
151
071
1;1
1@1
0B1
1c1
0e1
1i1
1n1
0p1
132
052
192
1>2
0@2
1a2
0c2
1g2
1l2
0n2
113
033
173
1<3
0>3
1_3
0a3
1e3
1j3
0l3
1/4
014
154
1:4
0<4
1]4
0_4
1c4
1h4
0j4
1-5
0/5
135
185
0:5
1[5
0]5
1a5
1f5
0h5
1+6
0-6
116
166
086
1Y6
0[6
1_6
1d6
0f6
1)7
0+7
1/7
147
067
1W7
0Y7
1]7
1b7
0d7
1'8
0)8
1-8
128
048
1U8
0W8
1[8
1`8
0b8
1%9
0'9
1+9
109
029
1S9
0U9
1Y9
1^9
0`9
1#:
0%:
1):
1.:
00:
1Q:
0S:
1W:
1\:
0^:
1!;
0#;
1';
1,;
0.;
1O;
0Q;
1U;
1Z;
0\;
1};
0!<
1%<
1*<
0,<
1M<
0O<
1S<
1X<
0Z<
1{<
0}<
1#=
1(=
0*=
1K=
0M=
1Q=
1V=
0X=
1y=
0{=
1!>
1&>
0(>
1I>
0K>
1O>
1T>
0V>
1w>
0y>
1}>
1$?
0&?
1G?
0I?
1M?
1R?
0T?
1u?
0w?
1{?
1"@
0$@
1E@
0G@
1K@
1P@
0R@
1I
0p
0@"
0n"
1E#
0l#
0<$
0j$
0:%
0h%
08&
0f&
06'
0d'
04(
0b(
02)
0`)
00*
0^*
0.+
0\+
0,,
0Z,
0*-
0X-
0(.
0V.
0&/
0T/
0$0
0R0
0"1
0P1
0~1
0N2
0|2
0L3
0z3
0J4
0x4
0H5
0v5
0F6
0t6
0D7
0r7
0B8
0p8
0@9
0n9
0>:
0l:
0<;
0j;
0:<
0h<
08=
0f=
06>
0d>
04?
0b?
02@
1E
0o
0?"
0m"
0=#
0k#
0;$
0i$
1=%
0g%
07&
0e&
05'
0c'
03(
0a(
01)
0_)
0/*
0]*
0-+
0[+
0+,
0Y,
0)-
0W-
0'.
0U.
0%/
0S/
0#0
0Q0
0!1
0O1
0}1
0M2
0{2
0K3
0y3
0I4
0w4
0G5
0u5
0E6
0s6
0C7
0q7
0A8
0o8
0?9
0m9
0=:
0k:
0;;
0i;
09<
0g<
07=
0e=
05>
0c>
03?
0a?
01@
0T
0Z
0_
0$"
0*"
0/"
0R"
0X"
0]"
0"#
0(#
0-#
0P#
0V#
0[#
0~#
0&$
0+$
0N$
0T$
0Y$
0|$
0$%
0)%
0L%
0R%
0W%
0z%
0"&
0'&
0J&
0P&
0U&
0x&
0~&
0%'
0H'
0N'
0S'
0v'
0|'
0#(
0F(
0L(
0Q(
0t(
0z(
0!)
0D)
0J)
0O)
0r)
0x)
0})
0B*
0H*
0M*
0p*
0v*
0{*
0@+
0F+
0K+
0n+
0t+
0y+
0>,
0D,
0I,
0l,
0r,
0w,
0<-
0B-
0G-
0j-
0p-
0u-
0:.
0@.
0E.
0h.
0n.
0s.
08/
0>/
0C/
0f/
0l/
0q/
060
0<0
0A0
0d0
0j0
0o0
041
0:1
0?1
0b1
0h1
0m1
022
082
0=2
0`2
0f2
0k2
003
063
0;3
0^3
0d3
0i3
0.4
044
094
0\4
0b4
0g4
0,5
025
075
0Z5
0`5
0e5
0*6
006
056
0X6
0^6
0c6
0(7
0.7
037
0V7
0\7
0a7
0&8
0,8
018
0T8
0Z8
0_8
0$9
0*9
0/9
0R9
0X9
0]9
0":
0(:
0-:
0P:
0V:
0[:
0~:
0&;
0+;
0N;
0T;
0Y;
0|;
0$<
0)<
0L<
0R<
0W<
0z<
0"=
0'=
0J=
0P=
0U=
0x=
0~=
0%>
0H>
0N>
0S>
0v>
0|>
0#?
0F?
0L?
0Q?
0t?
0z?
0!@
0D@
0J@
0O@
1H
0N
1v
0x
1F"
0H"
1t"
0v"
1D#
1r#
0t#
1B$
0D$
1p$
0r$
1@%
0B%
1n%
0p%
1>&
0@&
1l&
0n&
1<'
0>'
1j'
0l'
1:(
0<(
1h(
0j(
18)
0:)
1f)
0h)
16*
08*
1d*
0f*
14+
06+
1b+
0d+
12,
04,
1`,
0b,
10-
02-
1^-
0`-
1..
00.
1\.
0^.
1,/
0./
1Z/
0\/
1*0
0,0
1X0
0Z0
1(1
0*1
1V1
0X1
1&2
0(2
1T2
0V2
1$3
0&3
1R3
0T3
1"4
0$4
1P4
0R4
1~4
0"5
1N5
0P5
1|5
0~5
1L6
0N6
1z6
0|6
1J7
0L7
1x7
0z7
1H8
0J8
1v8
0x8
1F9
0H9
1t9
0v9
1D:
0F:
1r:
0t:
1B;
0D;
1p;
0r;
1@<
0B<
1n<
0p<
1>=
0@=
1l=
0n=
1<>
0>>
1j>
0l>
1:?
0<?
1h?
0j?
18@
0:@
1D
1r
0t
1B"
0D"
1p"
0r"
1@#
0B#
1n#
0p#
1>$
0@$
1l$
0n$
1<%
1j%
0l%
1:&
0<&
1h&
0j&
18'
0:'
1f'
0h'
16(
08(
1d(
0f(
14)
06)
1b)
0d)
12*
04*
1`*
0b*
10+
02+
1^+
0`+
1.,
00,
1\,
0^,
1,-
0.-
1Z-
0\-
1*.
0,.
1X.
0Z.
1(/
0*/
1V/
0X/
1&0
0(0
1T0
0V0
1$1
0&1
1R1
0T1
1"2
0$2
1P2
0R2
1~2
0"3
1N3
0P3
1|3
0~3
1L4
0N4
1z4
0|4
1J5
0L5
1x5
0z5
1H6
0J6
1v6
0x6
1F7
0H7
1t7
0v7
1D8
0F8
1r8
0t8
1B9
0D9
1p9
0r9
1@:
0B:
1n:
0p:
1>;
0@;
1l;
0n;
1<<
0><
1j<
0l<
1:=
0<=
1h=
0j=
18>
0:>
1f>
0h>
16?
08?
1d?
0f?
14@
06@
b0 :
b0 P
b0 h
b0 ~
b0 8"
b0 N"
b0 f"
b0 |"
b0 6#
b0 L#
b0 d#
b0 z#
b0 4$
b0 J$
b0 b$
b0 x$
b0 2%
b0 H%
b0 `%
b0 v%
b0 0&
b0 F&
b0 ^&
b0 t&
b0 .'
b0 D'
b0 \'
b0 r'
b0 ,(
b0 B(
b0 Z(
b0 p(
b0 *)
b0 @)
b0 X)
b0 n)
b0 (*
b0 >*
b0 V*
b0 l*
b0 &+
b0 <+
b0 T+
b0 j+
b0 $,
b0 :,
b0 R,
b0 h,
b0 "-
b0 8-
b0 P-
b0 f-
b0 ~-
b0 6.
b0 N.
b0 d.
b0 |.
b0 4/
b0 L/
b0 b/
b0 z/
b0 20
b0 J0
b0 `0
b0 x0
b0 01
b0 H1
b0 ^1
b0 v1
b0 .2
b0 F2
b0 \2
b0 t2
b0 ,3
b0 D3
b0 Z3
b0 r3
b0 *4
b0 B4
b0 X4
b0 p4
b0 (5
b0 @5
b0 V5
b0 n5
b0 &6
b0 >6
b0 T6
b0 l6
b0 $7
b0 <7
b0 R7
b0 j7
b0 "8
b0 :8
b0 P8
b0 h8
b0 ~8
b0 89
b0 N9
b0 f9
b0 |9
b0 6:
b0 L:
b0 d:
b0 z:
b0 4;
b0 J;
b0 b;
b0 x;
b0 2<
b0 H<
b0 `<
b0 v<
b0 0=
b0 F=
b0 ^=
b0 t=
b0 .>
b0 D>
b0 \>
b0 r>
b0 ,?
b0 B?
b0 Z?
b0 p?
b0 *@
b0 @@
07
08
0d
04"
0b"
02#
0`#
00$
0^$
0.%
0\%
0,&
0Z&
0*'
0X'
0((
0V(
0&)
0T)
0$*
0R*
0"+
0P+
0~+
0N,
0|,
0L-
0z-
0J.
0x.
0H/
0v/
0F0
0t0
0D1
0r1
0B2
0p2
0@3
0n3
0>4
0l4
0<5
0j5
0:6
0h6
087
0f7
068
0d8
049
0b9
02:
0`:
00;
0^;
0.<
0\<
0,=
0Z=
0*>
0X>
0(?
0V?
0&@
06
0c
03"
0a"
01#
0_#
0/$
0]$
0-%
0[%
0+&
0Y&
0)'
0W'
0'(
0U(
0%)
0S)
0#*
0Q*
0!+
0O+
0}+
0M,
0{,
0K-
0y-
0I.
0w.
0G/
0u/
0E0
0s0
0C1
0q1
0A2
0o2
0?3
0m3
0=4
0k4
0;5
0i5
096
0g6
077
0e7
058
0c8
039
0a9
01:
0_:
0/;
0];
0-<
0[<
0+=
0Y=
0)>
0W>
0'?
0U?
0%@
b0 !
b0 *
b0 0
b0 /
0J
0F#
0F
0>%
0w
0G"
0u"
0s#
0C$
0q$
0A%
0o%
0?&
0m&
0='
0k'
0;(
0i(
09)
0g)
07*
0e*
05+
0c+
03,
0a,
01-
0_-
0/.
0].
0-/
0[/
0+0
0Y0
0)1
0W1
0'2
0U2
0%3
0S3
0#4
0Q4
0!5
0O5
0}5
0M6
0{6
0K7
0y7
0I8
0w8
0G9
0u9
0E:
0s:
0C;
0q;
0A<
0o<
0?=
0m=
0=>
0k>
0;?
0i?
09@
0s
0C"
0q"
0A#
0o#
0?$
0m$
0k%
0;&
0i&
09'
0g'
07(
0e(
05)
0c)
03*
0a*
01+
0_+
0/,
0],
0--
0[-
0+.
0Y.
0)/
0W/
0'0
0U0
0%1
0S1
0#2
0Q2
0!3
0O3
0}3
0M4
0{4
0K5
0y5
0I6
0w6
0G7
0u7
0E8
0s8
0C9
0q9
0A:
0o:
0?;
0m;
0=<
0k<
0;=
0i=
09>
0g>
07?
0e?
05@
b1 ?
b1 G
1=
b10 m
b10 u
0k
b10 ="
b10 E"
0;"
b10 k"
b10 s"
0i"
b1 ;#
b1 C#
19#
b10 i#
b10 q#
0g#
b10 9$
b10 A$
07$
b10 g$
b10 o$
0e$
b10 7%
b10 ?%
05%
b10 e%
b10 m%
0c%
b10 5&
b10 =&
03&
b10 c&
b10 k&
0a&
b10 3'
b10 ;'
01'
b10 a'
b10 i'
0_'
b10 1(
b10 9(
0/(
b10 _(
b10 g(
0](
b10 /)
b10 7)
0-)
b10 ])
b10 e)
0[)
b10 -*
b10 5*
0+*
b10 [*
b10 c*
0Y*
b10 ++
b10 3+
0)+
b10 Y+
b10 a+
0W+
b10 ),
b10 1,
0',
b10 W,
b10 _,
0U,
b10 '-
b10 /-
0%-
b10 U-
b10 ]-
0S-
b10 %.
b10 -.
0#.
b10 S.
b10 [.
0Q.
b10 #/
b10 +/
0!/
b10 Q/
b10 Y/
0O/
b10 !0
b10 )0
0}/
b10 O0
b10 W0
0M0
b10 }0
b10 '1
0{0
b10 M1
b10 U1
0K1
b10 {1
b10 %2
0y1
b10 K2
b10 S2
0I2
b10 y2
b10 #3
0w2
b10 I3
b10 Q3
0G3
b10 w3
b10 !4
0u3
b10 G4
b10 O4
0E4
b10 u4
b10 }4
0s4
b10 E5
b10 M5
0C5
b10 s5
b10 {5
0q5
b10 C6
b10 K6
0A6
b10 q6
b10 y6
0o6
b10 A7
b10 I7
0?7
b10 o7
b10 w7
0m7
b10 ?8
b10 G8
0=8
b10 m8
b10 u8
0k8
b10 =9
b10 E9
0;9
b10 k9
b10 s9
0i9
b10 ;:
b10 C:
09:
b10 i:
b10 q:
0g:
b10 9;
b10 A;
07;
b10 g;
b10 o;
0e;
b10 7<
b10 ?<
05<
b10 e<
b10 m<
0c<
b10 5=
b10 ==
03=
b10 c=
b10 k=
0a=
b10 3>
b10 ;>
01>
b10 a>
b10 i>
0_>
b10 1?
b10 9?
0/?
b10 _?
b10 g?
0]?
b10 /@
b10 7@
0-@
b1 >
b1 C
1<
b10 l
b10 q
0j
b10 <"
b10 A"
0:"
b10 j"
b10 o"
0h"
b10 :#
b10 ?#
08#
b10 h#
b10 m#
0f#
b10 8$
b10 =$
06$
b10 f$
b10 k$
0d$
b1 6%
b1 ;%
14%
b10 d%
b10 i%
0b%
b10 4&
b10 9&
02&
b10 b&
b10 g&
0`&
b10 2'
b10 7'
00'
b10 `'
b10 e'
0^'
b10 0(
b10 5(
0.(
b10 ^(
b10 c(
0\(
b10 .)
b10 3)
0,)
b10 \)
b10 a)
0Z)
b10 ,*
b10 1*
0**
b10 Z*
b10 _*
0X*
b10 *+
b10 /+
0(+
b10 X+
b10 ]+
0V+
b10 (,
b10 -,
0&,
b10 V,
b10 [,
0T,
b10 &-
b10 +-
0$-
b10 T-
b10 Y-
0R-
b10 $.
b10 ).
0".
b10 R.
b10 W.
0P.
b10 "/
b10 '/
0~.
b10 P/
b10 U/
0N/
b10 ~/
b10 %0
0|/
b10 N0
b10 S0
0L0
b10 |0
b10 #1
0z0
b10 L1
b10 Q1
0J1
b10 z1
b10 !2
0x1
b10 J2
b10 O2
0H2
b10 x2
b10 }2
0v2
b10 H3
b10 M3
0F3
b10 v3
b10 {3
0t3
b10 F4
b10 K4
0D4
b10 t4
b10 y4
0r4
b10 D5
b10 I5
0B5
b10 r5
b10 w5
0p5
b10 B6
b10 G6
0@6
b10 p6
b10 u6
0n6
b10 @7
b10 E7
0>7
b10 n7
b10 s7
0l7
b10 >8
b10 C8
0<8
b10 l8
b10 q8
0j8
b10 <9
b10 A9
0:9
b10 j9
b10 o9
0h9
b10 ::
b10 ?:
08:
b10 h:
b10 m:
0f:
b10 8;
b10 =;
06;
b10 f;
b10 k;
0d;
b10 6<
b10 ;<
04<
b10 d<
b10 i<
0b<
b10 4=
b10 9=
02=
b10 b=
b10 g=
0`=
b10 2>
b10 7>
00>
b10 `>
b10 e>
0^>
b10 0?
b10 5?
0.?
b10 ^?
b10 c?
0\?
b10 .@
b10 3@
0,@
b11100 '
b11100 .
b11111 &
b11111 -
b10 %
b10 ,
b10011111000011100 +
b10001 )
b10001 5
b100000001 (
b100000001 4
#10
0;
0a
1/'
1]'
1-(
1[(
1+)
1Y)
1)*
1W*
1'+
1U+
1%,
1S,
1#-
1Q-
1!.
1O.
1}.
1M/
1{/
1K0
1y0
1I1
1w1
1G2
1u2
1E3
1s3
1C4
1q4
1A5
1o5
1?6
1m6
1=7
1k7
1;8
1i8
199
1g9
17:
1e:
15;
1c;
13<
1a<
11=
1_=
1/>
1]>
1-?
1[?
1Y
1+@
1U'
1%(
1S(
1#)
1Q)
1!*
1O*
1}*
1M+
1{+
1K,
1y,
1I-
1w-
1G.
1u.
1E/
1s/
1C0
1q0
1A1
1o1
1?2
1m2
1=3
1k3
1;4
1i4
195
1g5
176
1e6
157
1c7
138
1a8
119
1_9
1/:
1]:
1-;
1[;
1+<
1Y<
1)=
1W=
1'>
1U>
1%?
1S?
1#@
1]
1Q@
b0 ("
0S
b10 Q
b10 ^
0y
b1 z'
1G'
b1 J(
1u'
b1 s'
b1 "(
b1 x(
1E(
b1 C(
b1 P(
b1 H)
1s(
b1 q(
b1 ~(
b1 v)
1C)
b1 A)
b1 N)
b1 F*
1q)
b1 o)
b1 |)
b1 t*
1A*
b1 ?*
b1 L*
b1 D+
1o*
b1 m*
b1 z*
b1 r+
1?+
b1 =+
b1 J+
b1 B,
1m+
b1 k+
b1 x+
b1 p,
1=,
b1 ;,
b1 H,
b1 @-
1k,
b1 i,
b1 v,
b1 n-
1;-
b1 9-
b1 F-
b1 >.
1i-
b1 g-
b1 t-
b1 l.
b1 X8
19.
b1 7.
b1 D.
b1 </
b1 |=
1g.
b1 e.
b1 r.
b1 j/
17/
b1 5/
b1 B/
b1 :0
1e/
b1 c/
b1 p/
b1 h0
150
b1 30
b1 @0
b1 81
1c0
b1 a0
b1 n0
b1 f1
131
b1 11
b1 >1
b1 62
1a1
b1 _1
b1 l1
b1 d2
112
b1 /2
b1 <2
b1 43
1_2
b1 ]2
b1 j2
b1 b3
1/3
b1 -3
b1 :3
b1 24
1]3
b1 [3
b1 h3
b1 `4
1-4
b1 +4
b1 84
b1 05
1[4
b1 Y4
b1 f4
b1 ^5
1+5
b1 )5
b1 65
b1 .6
1Y5
b1 W5
b1 d5
b1 \6
1)6
b1 '6
b1 46
b1 ,7
1W6
b1 U6
b1 b6
b1 Z7
1'7
b1 %7
b1 27
b1 *8
1U7
b1 S7
b1 `7
1%8
b1 #8
b1 08
b1 (9
1S8
b1 Q8
b1 ^8
b1 V9
1#9
b1 !9
b1 .9
b1 &:
1Q9
b1 O9
b1 \9
b1 T:
1!:
b1 }9
b1 ,:
b1 $;
1O:
b1 M:
b1 Z:
b1 R;
1}:
b1 {:
b1 *;
b1 "<
1M;
b1 K;
b1 X;
b1 P<
1{;
b1 y;
b1 (<
b1 ~<
1K<
b1 I<
b1 V<
b1 N=
1y<
b1 w<
b1 &=
1I=
b1 G=
b1 T=
b1 L>
1w=
b1 u=
b1 $>
b1 z>
1G>
b1 E>
b1 R>
b1 J?
1u>
b1 s>
b1 "?
b1 x?
1E?
b1 C?
b1 P?
b1 H@
1s?
b1 q?
b1 ~?
1C@
b1 A@
b1 N@
17#
1e#
15$
1c$
13%
1a%
11&
1_&
0e
1m'
1K'
1=(
1y'
1k(
1I(
1;)
1w(
1i)
1G)
19*
1u)
1g*
1E*
17+
1s*
1e+
1C+
15,
1q+
1c,
1A,
13-
1o,
1a-
1?-
11.
1m-
1_.
1K8
1=.
1//
1o=
1k.
1]/
1;/
1-0
1i/
1[0
190
1+1
1g0
1Y1
171
1)2
1e1
1W2
152
1'3
1c2
1U3
133
1%4
1a3
1S4
114
1#5
1_4
1Q5
1/5
1!6
1]5
1O6
1-6
1}6
1[6
1M7
1+7
1{7
1Y7
1)8
1y8
1W8
1I9
1'9
1w9
1U9
1G:
1%:
1u:
1S:
1E;
1#;
1s;
1Q;
1C<
1!<
1q<
1O<
1A=
1}<
1M=
1?>
1{=
1m>
1K>
1=?
1y>
1k?
1I?
1;@
1w?
13
1G@
1]#
1-$
1[$
1+%
1Y%
1)&
1W&
1''
09
b0 R
1Y'
1)(
1W(
1')
1U)
1%*
1S*
1#+
1Q+
1!,
1O,
1},
1M-
1{-
1K.
178
1y.
1[=
1I/
1w/
1G0
1u0
1E1
1s1
1C2
1q2
1A3
1o3
1?4
1m4
1=5
1k5
1;6
1i6
197
1g7
1e8
159
1c9
13:
1a:
11;
1_;
1/<
1]<
1-=
1+>
1Y>
1)?
1W?
1'@
0"
0)"
0M
b10 N#
1,'
b11 F'
1Z'
b11 t'
1*(
b11 D(
1X(
b11 r(
1()
b11 B)
1V)
b11 p)
1&*
b11 @*
1T*
b11 n*
1$+
b11 >+
1R+
b11 l+
1",
b11 <,
1P,
b11 j,
1~,
b11 :-
1N-
b11 h-
1|-
b11 8.
1L.
b11 f.
1z.
b11 6/
1J/
b11 d/
1x/
b11 40
1H0
b11 b0
1v0
b11 21
1F1
b11 `1
1t1
b11 02
1D2
b11 ^2
1r2
b11 .3
1B3
b11 \3
1p3
b11 ,4
1@4
b11 Z4
1n4
b11 *5
1>5
b11 X5
1l5
b11 (6
1<6
b11 V6
1j6
b11 &7
1:7
b11 T7
1h7
b11 $8
188
b11 R8
1f8
b11 "9
169
b11 P9
1d9
b11 ~9
14:
b11 N:
1b:
b11 |:
12;
b11 L;
1`;
b11 z;
10<
b11 J<
1^<
b11 x<
1.=
b11 H=
1\=
b11 v=
1,>
b11 F>
1Z>
b11 t>
1*?
b11 D?
1X?
b11 r?
1(@
b11 B@
0V
0,"
1O#
1}#
1M$
1{$
1K%
1y%
1I&
1w&
0B
0>#
0A
1H#
0I#
0w#
0G$
0u$
09%
1A'
1o'
b111 b'
b111 q'
1?(
b111 2(
b111 A(
1m(
b111 `(
b111 o(
1=)
b111 0)
b111 ?)
1k)
b111 ^)
b111 m)
1;*
b111 .*
b111 =*
1i*
b111 \*
b111 k*
19+
b111 ,+
b111 ;+
1g+
b111 Z+
b111 i+
17,
b111 *,
b111 9,
1e,
b111 X,
b111 g,
15-
b111 (-
b111 7-
1c-
b111 V-
b111 e-
13.
b111 &.
b111 5.
1a.
b111 T.
b111 c.
11/
b111 $/
b111 3/
1_/
b111 R/
b111 a/
1/0
b111 "0
b111 10
1]0
b111 P0
b111 _0
1-1
b111 ~0
b111 /1
1[1
b111 N1
b111 ]1
1+2
b111 |1
b111 -2
1Y2
b111 L2
b111 [2
1)3
b111 z2
b111 +3
1W3
b111 J3
b111 Y3
1'4
b111 x3
b111 )4
1U4
b111 H4
b111 W4
1%5
b111 v4
b111 '5
1S5
b111 F5
b111 U5
1#6
b111 t5
b111 %6
1Q6
b111 D6
b111 S6
1!7
b111 r6
b111 #7
1O7
b111 B7
b111 Q7
1}7
b111 p7
b111 !8
1M8
b111 @8
b111 O8
1{8
b111 n8
b111 }8
1K9
b111 >9
b111 M9
1y9
b111 l9
b111 {9
1I:
b111 <:
b111 K:
1w:
b111 j:
b111 y:
1G;
b111 :;
b111 I;
1u;
b111 h;
b111 w;
1E<
b111 8<
b111 G<
1s<
b111 f<
b111 u<
1C=
b111 6=
b111 E=
1q=
b111 d=
b111 s=
1A>
b111 4>
b111 C>
1o>
b111 b>
b111 q>
1??
b111 2?
b111 A?
1m?
b111 `?
b111 o?
1=@
b111 0@
b111 ?@
0U
0W
0[
0%"
0'"
0+"
0S"
0U"
0Y"
0##
0%#
0)#
0Q#
1S#
0W#
0!$
1#$
0'$
0O$
1Q$
0U$
0}$
1!%
0%%
0M%
1O%
0S%
0{%
1}%
0#&
0K&
1M&
0Q&
0y&
1{&
0!'
0I'
0O'
0w'
0}'
0G(
0M(
0u(
0{(
0E)
0K)
0s)
0y)
0C*
0I*
0q*
0w*
0A+
0G+
0o+
0u+
0?,
0E,
0m,
0s,
0=-
0C-
0k-
0q-
0;.
0A.
0i.
0o.
09/
0?/
0g/
0m/
070
0=0
0e0
0k0
051
0;1
0c1
0i1
032
092
0a2
0g2
013
073
0_3
0e3
0/4
054
0]4
0c4
0-5
035
0[5
0a5
0+6
016
0Y6
0_6
0)7
0/7
0W7
0]7
0'8
0-8
0U8
0[8
0%9
0+9
0S9
0Y9
0#:
0):
0Q:
0W:
0!;
0';
0O;
0U;
0};
0%<
0M<
0S<
0{<
0#=
0K=
0Q=
0y=
0!>
0I>
0O>
0w>
0}>
0G?
0M?
0u?
0{?
0E@
0K@
0I
b11 X
0E#
1:%
1h%
18&
1f&
16'
1d'
14(
1b(
12)
1`)
10*
1^*
1.+
1\+
1,,
1Z,
1*-
1X-
1(.
1V.
1&/
1T/
1$0
1R0
1"1
1P1
1~1
1N2
1|2
1L3
1z3
1J4
1x4
1H5
1v5
1F6
1t6
1D7
1r7
1B8
1p8
1@9
1n9
1>:
1l:
1<;
1j;
1:<
1h<
18=
1f=
16>
1d>
14?
1b?
12@
0E
1=#
1k#
1;$
1i$
0=%
15'
1c'
13(
1a(
11)
1_)
1/*
1]*
1-+
1[+
1+,
1Y,
1)-
1W-
1'.
1U.
1%/
1S/
1#0
1Q0
1!1
1O1
1}1
1M2
1{2
1K3
1y3
1I4
1w4
1G5
1u5
1E6
1s6
1C7
1q7
1A8
1o8
1?9
1m9
1=:
1k:
1;;
1i;
19<
1g<
17=
1e=
15>
1c>
13?
1a?
11@
1T
1Z
1$"
1*"
1R"
1X"
1"#
1(#
1P#
1V#
1~#
1&$
1N$
1T$
1|$
1$%
1L%
1R%
1z%
1"&
1J&
1P&
1x&
1~&
1H'
1N'
1v'
1|'
1F(
1L(
1t(
1z(
1D)
1J)
1r)
1x)
1B*
1H*
1p*
1v*
1@+
1F+
1n+
1t+
1>,
1D,
1l,
1r,
1<-
1B-
1j-
1p-
1:.
1@.
1h.
1n.
18/
1>/
1f/
1l/
160
1<0
1d0
1j0
141
1:1
1b1
1h1
122
182
1`2
1f2
103
163
1^3
1d3
1.4
144
1\4
1b4
1,5
125
1Z5
1`5
1*6
106
1X6
1^6
1(7
1.7
1V7
1\7
1&8
1,8
1T8
1Z8
1$9
1*9
1R9
1X9
1":
1(:
1P:
1V:
1~:
1&;
1N;
1T;
1|;
1$<
1L<
1R<
1z<
1"=
1J=
1P=
1x=
1~=
1H>
1N>
1v>
1|>
1F?
1L?
1t?
1z?
1D@
1J@
0H
1K
b1100 @
b1100 O
0v
0F"
0t"
0D#
0r#
0B$
0p$
0@%
1B%
0n%
1p%
0>&
1@&
0l&
1n&
0<'
1>'
0j'
1l'
0:(
1<(
0h(
1j(
08)
1:)
0f)
1h)
06*
18*
0d*
1f*
04+
16+
0b+
1d+
02,
14,
0`,
1b,
00-
12-
0^-
1`-
0..
10.
0\.
1^.
0,/
1./
0Z/
1\/
0*0
1,0
0X0
1Z0
0(1
1*1
0V1
1X1
0&2
1(2
0T2
1V2
0$3
1&3
0R3
1T3
0"4
1$4
0P4
1R4
0~4
1"5
0N5
1P5
0|5
1~5
0L6
1N6
0z6
1|6
0J7
1L7
0x7
1z7
0H8
1J8
0v8
1x8
0F9
1H9
0t9
1v9
0D:
1F:
0r:
1t:
0B;
1D;
0p;
1r;
0@<
1B<
0n<
1p<
0>=
1@=
0l=
1n=
0<>
1>>
0j>
1l>
0:?
1<?
0h?
1j?
08@
1:@
0D
0r
0B"
0p"
0@#
1B#
0n#
1p#
0>$
1@$
0l$
1n$
0<%
0j%
0:&
0h&
08'
1:'
0f'
1h'
06(
18(
0d(
1f(
04)
16)
0b)
1d)
02*
14*
0`*
1b*
00+
12+
0^+
1`+
0.,
10,
0\,
1^,
0,-
1.-
0Z-
1\-
0*.
1,.
0X.
1Z.
0(/
1*/
0V/
1X/
0&0
1(0
0T0
1V0
0$1
1&1
0R1
1T1
0"2
1$2
0P2
1R2
0~2
1"3
0N3
1P3
0|3
1~3
0L4
1N4
0z4
1|4
0J5
1L5
0x5
1z5
0H6
1J6
0v6
1x6
0F7
1H7
0t7
1v7
0D8
1F8
0r8
1t8
0B9
1D9
0p9
1r9
0@:
1B:
0n:
1p:
0>;
1@;
0l;
1n;
0<<
1><
0j<
1l<
0:=
1<=
0h=
1j=
08>
1:>
0f>
1h>
06?
18?
0d?
1f?
04@
16@
b1 :
b1 P
b1 h
b1 ~
b1 8"
b1 N"
b1 f"
b1 |"
b1 6#
b1 L#
b1 d#
b1 z#
b1 4$
b1 J$
b1 b$
b1 x$
b1 2%
b1 H%
b1 `%
b1 v%
b1 0&
b1 F&
b1 ^&
b1 t&
b1 .'
b1 D'
b1 \'
b1 r'
b1 ,(
b1 B(
b1 Z(
b1 p(
b1 *)
b1 @)
b1 X)
b1 n)
b1 (*
b1 >*
b1 V*
b1 l*
b1 &+
b1 <+
b1 T+
b1 j+
b1 $,
b1 :,
b1 R,
b1 h,
b1 "-
b1 8-
b1 P-
b1 f-
b1 ~-
b1 6.
b1 N.
b1 d.
b1 |.
b1 4/
b1 L/
b1 b/
b1 z/
b1 20
b1 J0
b1 `0
b1 x0
b1 01
b1 H1
b1 ^1
b1 v1
b1 .2
b1 F2
b1 \2
b1 t2
b1 ,3
b1 D3
b1 Z3
b1 r3
b1 *4
b1 B4
b1 X4
b1 p4
b1 (5
b1 @5
b1 V5
b1 n5
b1 &6
b1 >6
b1 T6
b1 l6
b1 $7
b1 <7
b1 R7
b1 j7
b1 "8
b1 :8
b1 P8
b1 h8
b1 ~8
b1 89
b1 N9
b1 f9
b1 |9
b1 6:
b1 L:
b1 d:
b1 z:
b1 4;
b1 J;
b1 b;
b1 x;
b1 2<
b1 H<
b1 `<
b1 v<
b1 0=
b1 F=
b1 ^=
b1 t=
b1 .>
b1 D>
b1 \>
b1 r>
b1 ,?
b1 B?
b1 Z?
b1 p?
b1 *@
b1 @@
17
18
1d
14"
1b"
12#
1`#
10$
1^$
1.%
1\%
1,&
1Z&
1*'
1X'
1((
1V(
1&)
1T)
1$*
1R*
1"+
1P+
1~+
1N,
1|,
1L-
1z-
1J.
1x.
1H/
1v/
1F0
1t0
1D1
1r1
1B2
1p2
1@3
1n3
1>4
1l4
1<5
1j5
1:6
1h6
187
1f7
168
1d8
149
1b9
12:
1`:
10;
1^;
1.<
1\<
1,=
1Z=
1*>
1X>
1(?
1V?
1&@
16
1c
13"
1a"
11#
1_#
1/$
1]$
1-%
1[%
1+&
1Y&
1)'
1W'
1'(
1U(
1%)
1S)
1#*
1Q*
1!+
1O+
1}+
1M,
1{,
1K-
1y-
1I.
1w.
1G/
1u/
1E0
1s0
1C1
1q1
1A2
1o2
1?3
1m3
1=4
1k4
1;5
1i5
196
1g6
177
1e7
158
1c8
139
1a9
11:
1_:
1/;
1];
1-<
1[<
1+=
1Y=
1)>
1W>
1'?
1U?
1%@
b1101 !
b1101 *
b1101 0
b1101 /
0M'
b1 E'
b1 R'
0P'
b0 L'
0?'
b11 4'
b11 C'
0+'
0\&
0r&
0[&
0.&
0D&
0-&
0Q%
b1 I%
b1 V%
0^%
0T%
0t%
0]%
b1 P%
00%
1C%
b110 8%
b110 G%
0F%
0/%
0`$
0v$
0_$
02$
0H$
01$
0W"
0i
0'#
09"
0U#
b1 M#
b1 Z#
0b#
0g"
b1111111111111111111111111111111111111111111111111111111111110000 #
b1111111111111111111111111111111111111111111111111111111111110000 2
0Z"
01"
0*#
0_"
0X#
0x#
0/#
0%$
b1 {#
b1 *$
0S$
b1 K$
b1 X$
0#%
b1 y$
b1 (%
0a#
0!&
b1 w%
b1 &&
0O&
b1 G&
b1 T&
0}&
b1 u&
b1 $'
0($
0V$
0&%
b0 V"
0#"
b0 !"
b0 ."
b0 &#
0Q"
b0 O"
b0 \"
b1 T#
04#
0!#
b0 }"
b0 ,#
0$&
0R&
0"'
0I"
0&"
0w"
0T"
1G#
b110 <#
b110 K#
0J#
0$#
b1 $$
b1 R$
b1 "%
05"
0c"
03#
b1 ~%
b1 N&
b1 |&
1u#
b10 |#
1E$
b10 L$
1s$
b10 z$
0f
b0 ""
06"
b0 P"
0d"
b1111111111111111111111111111111111111111111111111111000000000000 1
b0 ~"
1q%
b10 x%
1A&
b10 H&
1o&
b10 v&
1v#
b110 j#
b110 y#
1F$
b110 :$
b110 I$
1t$
b110 h$
b110 w$
0{
b0 n
b0 }
0K"
b0 >"
b0 M"
0y"
b0 l"
b0 {"
1r%
b110 f%
b110 u%
1B&
b110 6&
b110 E&
1p&
b110 d&
b110 s&
0p
0@"
0n"
0l#
0<$
0j$
0o
0?"
0m"
0g%
07&
0e&
0w
0G"
0u"
0s#
0C$
0q$
0s
0C"
0q"
0k%
0;&
0i&
b1 m
b1 u
1k
b1 ="
b1 E"
1;"
b1 k"
b1 s"
1i"
b1 i#
b1 q#
1g#
b1 9$
b1 A$
17$
b1 g$
b1 o$
1e$
b1 l
b1 q
1j
b1 <"
b1 A"
1:"
b1 j"
b1 o"
1h"
b1 d%
b1 i%
1b%
b1 4&
b1 9&
12&
b1 b&
b1 g&
1`&
b111011100 '
b111011100 .
b10011111111011100 +
b11111111 )
b11111111 5
b111100001111 (
b111100001111 4
#15
1$
07#
0e#
05$
0c$
03%
0a%
01&
0_&
0/'
0]'
0-(
0[(
0+)
0Y)
0)*
0W*
0'+
0U+
0%,
0S,
0#-
0Q-
0!.
0O.
0}.
0M/
0{/
0K0
0y0
0I1
0w1
0G2
0u2
0E3
0s3
0C4
0q4
0A5
0o5
0?6
0m6
0=7
0k7
0;8
0i8
099
0g9
07:
05;
0c;
03<
1a<
01=
0_=
0/>
0-?
0[?
0Y
0+@
0]#
0-$
0[$
0+%
0Y%
0)&
0W&
0''
0U'
0%(
0S(
0#)
0Q)
0!*
0O*
0}*
0M+
0{+
0K,
0y,
0I-
0w-
0G.
0u.
0E/
0s/
0C0
0q0
0A1
0o1
0?2
0m2
0=3
0k3
0;4
0i4
095
0g5
076
0e6
057
0c7
038
0a8
019
0_9
0/:
0]:
0[;
0+<
0Y<
1)=
0W=
0'>
0U>
0S?
0#@
0]
0Q@
0O#
b0 M#
b0 Z#
0}#
b0 {#
b0 *$
0M$
b0 K$
b0 X$
0{$
b0 y$
b0 (%
0K%
b0 I%
b0 V%
0y%
b0 w%
b0 &&
0I&
b0 G&
b0 T&
0w&
b0 u&
b0 $'
b0 z'
0G'
b0 E'
b0 R'
b0 J(
0u'
b0 s'
b0 "(
b0 x(
0E(
b0 C(
b0 P(
b0 H)
0s(
b0 q(
b0 ~(
b0 v)
0C)
b0 A)
b0 N)
b0 F*
0q)
b0 o)
b0 |)
b0 t*
0A*
b0 ?*
b0 L*
b0 D+
0o*
b0 m*
b0 z*
b0 r+
0?+
b0 =+
b0 J+
b0 B,
0m+
b0 k+
b0 x+
b0 p,
0=,
b0 ;,
b0 H,
b0 @-
0k,
b0 i,
b0 v,
b0 n-
0;-
b0 9-
b0 F-
b0 >.
0i-
b0 g-
b0 t-
b0 l.
b0 X8
09.
b0 7.
b0 D.
b0 </
b0 |=
0g.
b0 e.
b0 r.
b0 j/
07/
b0 5/
b0 B/
b0 :0
0e/
b0 c/
b0 p/
b0 h0
050
b0 30
b0 @0
b0 81
0c0
b0 a0
b0 n0
b0 f1
031
b0 11
b0 >1
b0 62
0a1
b0 _1
b0 l1
b0 d2
012
b0 /2
b0 <2
b0 43
0_2
b0 ]2
b0 j2
b0 b3
0/3
b0 -3
b0 :3
b0 24
0]3
b0 [3
b0 h3
b0 `4
0-4
b0 +4
b0 84
b0 05
0[4
b0 Y4
b0 f4
b0 ^5
0+5
b0 )5
b0 65
b0 .6
0Y5
b0 W5
b0 d5
b0 \6
0)6
b0 '6
b0 46
b0 ,7
0W6
b0 U6
b0 b6
b0 Z7
0'7
b0 %7
b0 27
b0 *8
0U7
b0 S7
b0 `7
0%8
b0 #8
b0 08
b0 (9
0S8
b0 Q8
b0 ^8
b0 V9
0#9
b0 !9
b0 .9
b0 &:
0Q9
b0 O9
b0 \9
b0 T:
0!:
b0 }9
b0 ,:
0O:
b0 M:
b0 Z:
b0 "<
0M;
b0 K;
b0 X;
b0 P<
0{;
b0 y;
b0 (<
0K<
b0 I<
b0 V<
1y<
b1 w<
b1 &=
0I=
b0 G=
b0 T=
b0 L>
0w=
b0 u=
b0 $>
b0 z>
0G>
b0 E>
b0 R>
b0 x?
0E?
b0 C?
b0 P?
b0 H@
0s?
b0 q?
b0 ~?
0C@
b0 A@
b0 N@
0S#
0#$
0Q$
0!%
0O%
0}%
0M&
0{&
0m'
0K'
0=(
0y'
0k(
0I(
0;)
0w(
0i)
0G)
09*
0u)
0g*
0E*
07+
0s*
0e+
0C+
05,
0q+
0c,
0A,
03-
0o,
0a-
0?-
01.
0m-
0_.
0K8
0=.
0//
0o=
0k.
0]/
0;/
0-0
0i/
0[0
090
0+1
0g0
0Y1
071
0)2
0e1
0W2
052
0'3
0c2
0U3
033
0%4
0a3
0S4
014
0#5
0_4
0Q5
0/5
0!6
0]5
0O6
0-6
0}6
0[6
0M7
0+7
0{7
0Y7
0)8
0y8
0W8
0I9
0'9
0w9
0U9
0G:
0%:
0S:
0s;
0Q;
0C<
0!<
0O<
1}<
0M=
0?>
0{=
0m>
0K>
0k?
0I?
0;@
0w?
03
0G@
0Y'
0)(
0W(
0')
0U)
0%*
0S*
0#+
0Q+
0!,
0O,
0},
0M-
0{-
0K.
078
0y.
0[=
0I/
0w/
0G0
0u0
0E1
0s1
0C2
0q2
0A3
0o3
0?4
0m4
0=5
0k5
0;6
0i6
097
0g7
0e8
059
0c9
03:
0a:
0_;
0/<
0]<
0+>
0Y>
0W?
0'@
0"
0,'
b0 F'
0Z'
b0 t'
0*(
b0 D(
0X(
b0 r(
0()
b0 B)
0V)
b0 p)
0&*
b0 @*
0T*
b0 n*
0$+
b0 >+
0R+
b0 l+
0",
b0 <,
0P,
b0 j,
0~,
b0 :-
0N-
b0 h-
0|-
b0 8.
0L.
b0 f.
0z.
b0 6/
0J/
b0 d/
0x/
b0 40
0H0
b0 b0
0v0
b0 21
0F1
b0 `1
0t1
b0 02
0D2
b0 ^2
0r2
b0 .3
0B3
b0 \3
0p3
b0 ,4
0@4
b0 Z4
0n4
b0 *5
0>5
b0 X5
0l5
b0 (6
0<6
b0 V6
0j6
b0 &7
0:7
b0 T7
0h7
b0 $8
088
b0 R8
0f8
b0 "9
069
b0 P9
0d9
b0 ~9
04:
b0 N:
02;
b0 L;
0`;
b0 z;
00<
b0 J<
0.=
b0 H=
0\=
b0 v=
0,>
b0 F>
0*?
b0 D?
0X?
b0 r?
0(@
b0 B@
0A'
0o'
b0 b'
b0 q'
0?(
b0 2(
b0 A(
0m(
b0 `(
b0 o(
0=)
b0 0)
b0 ?)
0k)
b0 ^)
b0 m)
0;*
b0 .*
b0 =*
0i*
b0 \*
b0 k*
09+
b0 ,+
b0 ;+
0g+
b0 Z+
b0 i+
07,
b0 *,
b0 9,
0e,
b0 X,
b0 g,
05-
b0 (-
b0 7-
0c-
b0 V-
b0 e-
03.
b0 &.
b0 5.
0a.
b0 T.
b0 c.
01/
b0 $/
b0 3/
0_/
b0 R/
b0 a/
0/0
b0 "0
b0 10
0]0
b0 P0
b0 _0
0-1
b0 ~0
b0 /1
0[1
b0 N1
b0 ]1
0+2
b0 |1
b0 -2
0Y2
b0 L2
b0 [2
0)3
b0 z2
b0 +3
0W3
b0 J3
b0 Y3
0'4
b0 x3
b0 )4
0U4
b0 H4
b0 W4
0%5
b0 v4
b0 '5
0S5
b0 F5
b0 U5
0#6
b0 t5
b0 %6
0Q6
b0 D6
b0 S6
0!7
b0 r6
b0 #7
0O7
b0 B7
b0 Q7
0}7
b0 p7
b0 !8
0M8
b0 @8
b0 O8
0{8
b0 n8
b0 }8
0K9
b0 >9
b0 M9
0y9
b0 l9
b0 {9
0I:
b0 <:
b0 K:
0G;
0u;
b0 h;
b0 w;
0E<
b0 8<
b0 G<
0C=
0q=
b0 d=
b0 s=
0A>
b0 4>
b0 C>
0??
0m?
b0 `?
b0 o?
0=@
b0 0@
b0 ?@
b0 X
0:%
0h%
08&
0f&
06'
0d'
04(
0b(
02)
0`)
00*
0^*
0.+
0\+
0,,
0Z,
0*-
0X-
0(.
0V.
0&/
0T/
0$0
0R0
0"1
0P1
0~1
0N2
0|2
0L3
0z3
0J4
0x4
0H5
0v5
0F6
0t6
0D7
0r7
0B8
0p8
0@9
0n9
0>:
0l:
0<;
0j;
0:<
1o<
08=
0f=
06>
1k>
04?
0b?
02@
0=#
0k#
0;$
0i$
05'
0c'
03(
0a(
01)
0_)
0/*
0]*
0-+
0[+
0+,
0Y,
0)-
0W-
0'.
0U.
0%/
0S/
0#0
0Q0
0!1
0O1
0}1
0M2
0{2
0K3
0y3
0I4
0w4
0G5
0u5
0E6
0s6
0C7
0q7
0A8
0o8
0?9
0m9
0=:
1o:
0;;
0i;
09<
0g<
07=
0e=
05>
1g>
03?
0a?
01@
1H
0K
1v
1F"
1t"
1D#
1r#
1B$
1p$
1@%
0B%
1n%
0p%
1>&
0@&
1l&
0n&
1<'
0>'
1j'
0l'
1:(
0<(
1h(
0j(
18)
0:)
1f)
0h)
16*
08*
1d*
0f*
14+
06+
1b+
0d+
12,
04,
1`,
0b,
10-
02-
1^-
0`-
1..
00.
1\.
0^.
1,/
0./
1Z/
0\/
1*0
0,0
1X0
0Z0
1(1
0*1
1V1
0X1
1&2
0(2
1T2
0V2
1$3
0&3
1R3
0T3
1"4
0$4
1P4
0R4
1~4
0"5
1N5
0P5
1|5
0~5
1L6
0N6
1z6
0|6
1J7
0L7
1x7
0z7
1H8
0J8
1v8
0x8
1F9
0H9
1t9
0v9
1D:
0F:
1r:
0t:
1B;
0D;
1p;
0r;
1@<
0B<
1n<
1>=
0@=
1l=
0n=
1<>
0>>
1j>
1:?
0<?
1h?
0j?
18@
0:@
1D
1r
1B"
1p"
1@#
0B#
1n#
0p#
1>$
0@$
1l$
0n$
1<%
1j%
1:&
1h&
18'
0:'
1f'
0h'
16(
08(
1d(
0f(
14)
06)
1b)
0d)
12*
04*
1`*
0b*
10+
02+
1^+
0`+
1.,
00,
1\,
0^,
1,-
0.-
1Z-
0\-
1*.
0,.
1X.
0Z.
1(/
0*/
1V/
0X/
1&0
0(0
1T0
0V0
1$1
0&1
1R1
0T1
1"2
0$2
1P2
0R2
1~2
0"3
1N3
0P3
1|3
0~3
1L4
0N4
1z4
0|4
1J5
0L5
1x5
0z5
1H6
0J6
1v6
0x6
1F7
0H7
1t7
0v7
1D8
0F8
1r8
0t8
1B9
0D9
1p9
0r9
1@:
0B:
1n:
1>;
0@;
1l;
0n;
1<<
0><
1j<
0l<
1:=
0<=
1h=
0j=
18>
0:>
1f>
16?
08?
1d?
0f?
14@
06@
07
08
0d
04"
0b"
02#
0`#
00$
0^$
0.%
0\%
0,&
0Z&
0*'
0X'
0((
0V(
0&)
0T)
0$*
0R*
0"+
0P+
0~+
0N,
0|,
0L-
0z-
0J.
0x.
0H/
0v/
0F0
0t0
0D1
0r1
0B2
0p2
0@3
0n3
0>4
0l4
0<5
0j5
0:6
0h6
087
0f7
068
0d8
049
0b9
02:
0`:
00;
0^;
0.<
0\<
0,=
0Z=
0*>
0X>
0(?
0V?
0&@
06
0c
03"
0a"
01#
0_#
0/$
0]$
0-%
0[%
0+&
0Y&
0)'
0W'
0'(
0U(
0%)
0S)
0#*
0Q*
0!+
0O+
0}+
0M,
0{,
0K-
0y-
0I.
0w.
0G/
0u/
0E0
0s0
0C1
0q1
0A2
0o2
0?3
0m3
0=4
0k4
0;5
0i5
096
0g6
077
0e7
058
0c8
039
0a9
01:
0_:
0/;
0];
0-<
0[<
0+=
0Y=
0)>
0W>
0'?
0U?
0%@
b1 !
b1 *
b1 0
b1 /
0;
0i
09"
0g"
1]>
b1000100010000000000000000000000000000000000000000000000000000 #
b1000100010000000000000000000000000000000000000000000000000000 2
0a
01"
0_"
0/#
1%?
b0 N=
b0 ("
0S
b0 Q
b0 ^
b0 V"
0#"
b0 !"
b0 ."
b0 &#
0Q"
b0 O"
b0 \"
0!#
b0 }"
b0 ,#
b0 L'
b0 R;
b1 J?
1u>
b1 s>
b1 "?
0A=
b0 6=
b0 E=
0y
0W
0I"
0'"
0w"
0U"
0%#
0?'
b0 4'
b0 C'
0E;
b0 :;
b0 I;
1=?
b100 2?
b100 A?
1y>
b0 T#
0a#
b0 $$
01$
b0 R$
0_$
b0 "%
0/%
b1 ~<
0-=
0e
05"
0c"
03#
b0 P%
0]%
b0 ~%
0-&
b0 N&
0[&
b0 |&
0+'
b1 $;
01;
1)?
0G#
04#
b0 N#
0u#
0b#
b0 |#
0E$
02$
b0 L$
0s$
0`$
b0 z$
1q<
0t<
0^<
b10 x<
09
b0 R
0f
b0 ""
06"
b0 P"
0d"
b0 ~"
0C%
00%
b0 J%
0q%
0^%
b0 x%
0A&
0.&
b0 H&
0o&
0\&
b0 v&
1u:
0x:
0b:
b10 |:
1Z>
b1000000000000000000000000000000000000000000000000000000000000 1
b11 t>
0H#
0I#
b0 <#
b0 K#
0v#
0w#
b0 j#
b0 y#
0F$
0G$
b0 :$
b0 I$
0t$
0u$
b0 h$
b0 w$
1r<
0s<
b110 f<
b110 u<
0M
b0 @
b0 O
0{
b0 n
b0 }
0K"
b0 >"
b0 M"
0y"
b0 l"
b0 {"
0D%
0E%
b0 8%
b0 G%
0r%
0s%
b0 f%
b0 u%
0B&
0C&
b0 6&
b0 E&
0p&
0q&
b0 d&
b0 s&
1v:
0w:
b110 j:
b110 y:
1o>
b11 b>
b11 q>
0B
0p
0@"
0n"
0>#
0l#
0<$
0j$
1h<
1d>
0A
0o
0?"
0m"
09%
0g%
07&
0e&
1k:
1c>
0J
0x
0H"
0v"
0F#
0t#
0D$
0r$
0p<
0l>
0F
0t
0D"
0r"
0>%
0l%
0<&
0j&
0p:
0h>
b10 ?
b10 G
0=
b10 m
b10 u
0k
b10 ="
b10 E"
0;"
b10 k"
b10 s"
0i"
b10 ;#
b10 C#
09#
b10 i#
b10 q#
0g#
b10 9$
b10 A$
07$
b10 g$
b10 o$
0e$
b1 e<
b1 m<
1c<
b1 a>
b1 i>
1_>
b10 >
b10 C
0<
b10 l
b10 q
0j
b10 <"
b10 A"
0:"
b10 j"
b10 o"
0h"
b10 6%
b10 ;%
04%
b10 d%
b10 i%
0b%
b10 4&
b10 9&
02&
b10 b&
b10 g&
0`&
b1 h:
b1 m:
1f:
b1 `>
b1 e>
1^>
b110111100 '
b110111100 .
b10011111110111100 +
b1000100000000000000000000000000000000000000000000000000000000 )
b1000100000000000000000000000000000000000000000000000000000000 5
b1000000010000000000000000000000000000000000000000000000000000 (
b1000000010000000000000000000000000000000000000000000000000000 4
#20
1b
12"
10#
1Y
1)"
1'#
1\
1,"
1*#
1U
1[
0`
1%"
1+"
00"
1S"
1Y"
0^"
1##
1)#
0.#
1Q#
1W#
0\#
1!$
1'$
0,$
1O$
1U$
0Z$
1}$
1%%
0*%
1M%
1S%
0X%
1{%
1#&
0(&
1K&
1Q&
0V&
1y&
1!'
0&'
1I'
1O'
0T'
1w'
1}'
0$(
1G(
1M(
0R(
1u(
1{(
0")
1E)
1K)
0P)
1s)
1y)
0~)
1C*
1I*
0N*
1q*
1w*
0|*
1A+
1G+
0L+
1o+
1u+
0z+
1?,
1E,
0J,
1m,
1s,
0x,
1=-
1C-
0H-
1k-
1q-
0v-
1;.
1A.
0F.
1i.
1o.
0t.
19/
1?/
0D/
1g/
1m/
0r/
170
1=0
0B0
1e0
1k0
0p0
151
1;1
0@1
1c1
1i1
0n1
132
192
0>2
1a2
1g2
0l2
113
173
0<3
1_3
1e3
0j3
1/4
154
0:4
1]4
1c4
0h4
1-5
135
085
1[5
1a5
0f5
1+6
116
066
1Y6
1_6
0d6
1)7
1/7
047
1W7
1]7
0b7
1'8
1-8
028
1U8
1[8
0`8
1%9
1+9
009
1S9
1Y9
0^9
1#:
1):
0.:
1Q:
1W:
0\:
1!;
1';
0,;
1O;
1U;
0Z;
1};
1%<
0*<
1M<
1S<
0X<
1{<
1#=
0(=
1K=
1Q=
0V=
1y=
1!>
0&>
1I>
1O>
0T>
1w>
1}>
0$?
1G?
1M?
0R?
1u?
1{?
0"@
1E@
1K@
0P@
0T
0Z
1_
0$"
0*"
1/"
0R"
0X"
1]"
0"#
0(#
1-#
0P#
0V#
1[#
0~#
0&$
1+$
0N$
0T$
1Y$
0|$
0$%
1)%
0L%
0R%
1W%
0z%
0"&
1'&
0J&
0P&
1U&
0x&
0~&
1%'
0H'
0N'
1S'
0v'
0|'
1#(
0F(
0L(
1Q(
0t(
0z(
1!)
0D)
0J)
1O)
0r)
0x)
1})
0B*
0H*
1M*
0p*
0v*
1{*
0@+
0F+
1K+
0n+
0t+
1y+
0>,
0D,
1I,
0l,
0r,
1w,
0<-
0B-
1G-
0j-
0p-
1u-
0:.
0@.
1E.
0h.
0n.
1s.
08/
0>/
1C/
0f/
0l/
1q/
060
0<0
1A0
0d0
0j0
1o0
041
0:1
1?1
0b1
0h1
1m1
022
082
1=2
0`2
0f2
1k2
003
063
1;3
0^3
0d3
1i3
0.4
044
194
0\4
0b4
1g4
0,5
025
175
0Z5
0`5
1e5
0*6
006
156
0X6
0^6
1c6
0(7
0.7
137
0V7
0\7
1a7
0&8
0,8
118
0T8
0Z8
1_8
0$9
0*9
1/9
0R9
0X9
1]9
0":
0(:
1-:
0P:
0V:
1[:
0~:
0&;
1+;
0N;
0T;
1Y;
0|;
0$<
1)<
0L<
0R<
1W<
0z<
0"=
1'=
0J=
0P=
1U=
0x=
0~=
1%>
0H>
0N>
1S>
0v>
0|>
1#?
0F?
0L?
1Q?
0t?
0z?
1!@
0D@
0J@
1O@
b10 :
b10 P
b10 h
b10 ~
b10 8"
b10 N"
b10 f"
b10 |"
b10 6#
b10 L#
b10 d#
b10 z#
b10 4$
b10 J$
b10 b$
b10 x$
b10 2%
b10 H%
b10 `%
b10 v%
b10 0&
b10 F&
b10 ^&
b10 t&
b10 .'
b10 D'
b10 \'
b10 r'
b10 ,(
b10 B(
b10 Z(
b10 p(
b10 *)
b10 @)
b10 X)
b10 n)
b10 (*
b10 >*
b10 V*
b10 l*
b10 &+
b10 <+
b10 T+
b10 j+
b10 $,
b10 :,
b10 R,
b10 h,
b10 "-
b10 8-
b10 P-
b10 f-
b10 ~-
b10 6.
b10 N.
b10 d.
b10 |.
b10 4/
b10 L/
b10 b/
b10 z/
b10 20
b10 J0
b10 `0
b10 x0
b10 01
b10 H1
b10 ^1
b10 v1
b10 .2
b10 F2
b10 \2
b10 t2
b10 ,3
b10 D3
b10 Z3
b10 r3
b10 *4
b10 B4
b10 X4
b10 p4
b10 (5
b10 @5
b10 V5
b10 n5
b10 &6
b10 >6
b10 T6
b10 l6
b10 $7
b10 <7
b10 R7
b10 j7
b10 "8
b10 :8
b10 P8
b10 h8
b10 ~8
b10 89
b10 N9
b10 f9
b10 |9
b10 6:
b10 L:
b10 d:
b10 z:
b10 4;
b10 J;
b10 b;
b10 x;
b10 2<
b10 H<
b10 `<
b10 v<
b10 0=
b10 F=
b10 ^=
b10 t=
b10 .>
b10 D>
b10 \>
b10 r>
b10 ,?
b10 B?
b10 Z?
b10 p?
b10 *@
b10 @@
b10 !
b10 *
b10 0
b10 /
0$
1;
0a<
1i
1g"
0e:
0]>
b1011 #
b1011 2
0a
0)=
01"
0/#
0-;
0%?
0S
b10 Q
b10 ^
0y<
b0 w<
b0 &=
0#"
b10 !"
b10 ."
0!#
b10 }"
b10 ,#
0}:
b0 {:
b0 *;
b0 J?
0u>
b0 s>
b0 "?
0W
0}<
0'"
0%#
0#;
0=?
b0 2?
b0 A?
0y>
b1 X
b0 ~<
b1 ("
b1 &#
b0 $;
0)?
1K
b10 R
0q<
b0 x<
1y
b10 ""
1w"
b10 ~"
0u:
b0 |:
0Z>
b0 1
b0 t>
1L
b110 @
b110 O
0r<
b0 f<
b0 u<
1z
b110 n
b110 }
1x"
b110 l"
b110 {"
0v:
b0 j:
b0 y:
0o>
b0 b>
b0 q>
1B
0h<
0d>
1o
1m"
0k:
0c>
1I
0o<
0k>
1s
1q"
0o:
0g>
b1 ?
b1 G
1=
b10 e<
b10 m<
0c<
b10 a>
b10 i>
0_>
b1 l
b1 q
1j
b1 j"
b1 o"
1h"
b10 h:
b10 m:
0f:
b10 `>
b10 e>
0^>
b100001010 '
b100001010 .
b10011111100001010 +
b1 )
b1 5
b1010 (
b1010 4
#25
1h7
1~7
1g7
1:7
1P7
197
1j6
1"7
1i6
1<6
1R6
1;6
1l5
1$6
1k5
1>5
1T5
1=5
1n4
1&5
1m4
1@4
1V4
1?4
1p3
1(4
1o3
1B3
1.=
1X3
1D=
1A3
1-=
1r2
1^<
1*3
1t<
1q2
1]<
1D2
10<
1Z2
1F<
1C2
1/<
1t1
1`;
1,2
1v;
1s1
1_;
1F1
1(@
12;
1\1
0"
1>@
1H;
1E1
1'@
11;
1v0
1X?
1b:
1.1
1n?
1x:
1u0
1W?
1a:
1H0
1*?
14:
1^0
1@?
1J:
1G0
1)?
13:
1x/
1Z>
1d9
100
1p>
1z9
1w/
1Y>
1c9
1J/
1,>
169
1`/
1B>
1L9
1I/
1+>
159
1z.
1\=
1f8
12/
1r=
1|8
1y.
1[=
1e8
1L.
188
1b.
1N8
1K.
178
1|-
14.
1{-
1N-
1d-
1M-
1~,
16-
1},
1P,
1f,
1O,
1",
18,
1!,
1R+
1h+
1Q+
1$+
1:+
1#+
1T*
1j*
1S*
1&*
1<*
1%*
1V)
1l)
1U)
1()
1>)
1')
1X(
1n(
1W(
1*(
1@(
1)(
1Z'
1p'
1Y'
1,'
1B'
1+'
1\&
1r&
1[&
1.&
1D&
1-&
1^%
1t%
1]%
10%
1F%
1/%
1`$
1v$
1_$
12$
1H$
11$
1b#
07#
0e#
05$
0c$
03%
0a%
01&
0_&
0/'
0]'
0-(
0[(
0+)
0Y)
0)*
0W*
0'+
0U+
0%,
0S,
0#-
0Q-
0!.
0O.
0}.
0M/
0{/
0K0
0y0
0I1
0w1
0G2
0u2
0E3
0s3
0C4
0q4
0A5
0o5
0?6
0m6
0=7
0k7
0;8
0i8
099
0g9
07:
0e:
05;
0c;
03<
0a<
01=
0_=
0/>
0]>
0-?
0[?
0+@
1x#
0^#
0.$
0\$
0,%
0Z%
0*&
0X&
0('
0V'
0&(
0T(
0$)
0R)
0"*
0P*
0~*
0N+
0|+
0L,
0z,
0J-
0x-
0H.
0v.
0F/
0t/
0D0
0r0
0B1
0p1
0@2
0n2
0>3
0l3
0<4
0j4
0:5
0h5
086
0f6
067
0d7
048
0b8
029
0`9
00:
0^:
0.;
0\;
0,<
0Z<
0*=
0X=
0(>
0V>
0&?
0T?
0$@
0R@
1a#
14#
0U#
b0 M#
b0 Z#
0%$
b0 {#
b0 *$
0S$
b0 K$
b0 X$
0#%
b0 y$
b0 (%
0Q%
b0 I%
b0 V%
0!&
b0 w%
b0 &&
0O&
b0 G&
b0 T&
0}&
b0 u&
b0 $'
0M'
b0 E'
b0 R'
0{'
b0 s'
b0 "(
0K(
b0 C(
b0 P(
0y(
b0 q(
b0 ~(
0I)
b0 A)
b0 N)
0w)
b0 o)
b0 |)
0G*
b0 ?*
b0 L*
0u*
b0 m*
b0 z*
0E+
b0 =+
b0 J+
0s+
b0 k+
b0 x+
0C,
b0 ;,
b0 H,
0q,
b0 i,
b0 v,
0A-
b0 9-
b0 F-
0o-
b0 g-
b0 t-
0?.
b0 7.
b0 D.
0m.
b0 e.
b0 r.
0=/
b0 5/
b0 B/
0k/
b0 c/
b0 p/
0;0
b0 30
b0 @0
0i0
b0 a0
b0 n0
091
b0 11
b0 >1
0g1
b0 _1
b0 l1
072
b0 /2
b0 <2
0e2
b0 ]2
b0 j2
053
b0 -3
b0 :3
0c3
b0 [3
b0 h3
034
b0 +4
b0 84
0a4
b0 Y4
b0 f4
015
b0 )5
b0 65
0_5
b0 W5
b0 d5
0/6
b0 '6
b0 46
0]6
b0 U6
b0 b6
0-7
b0 %7
b0 27
0[7
b0 S7
b0 `7
0+8
b0 #8
b0 08
0Y8
b0 Q8
b0 ^8
0)9
b0 !9
b0 .9
0W9
b0 O9
b0 \9
0':
b0 }9
b0 ,:
0U:
b0 M:
b0 Z:
0%;
b0 {:
b0 *;
0S;
b0 K;
b0 X;
0#<
b0 y;
b0 (<
0Q<
b0 I<
b0 V<
0!=
b0 w<
b0 &=
0O=
b0 G=
b0 T=
0}=
b0 u=
b0 $>
0M>
b0 E>
b0 R>
0{>
b0 s>
b0 "?
0K?
b0 C?
b0 P?
0y?
b0 q?
b0 ~?
0I@
b0 A@
b0 N@
1#"
1Q"
1J#
0X#
0($
0V$
0&%
0T%
0$&
0R&
0"'
0P'
0~'
0N(
0|(
0L)
0z)
0J*
0x*
0H+
0v+
0F,
0t,
0D-
0r-
0B.
0p.
0@/
0n/
0>0
0l0
0<1
0j1
0:2
0h2
083
0f3
064
0d4
045
0b5
026
0`6
007
0^7
0.8
0\8
0,9
0Z9
0*:
0X:
0(;
0V;
0&<
0T<
0$=
0R=
0">
0P>
0~>
0N?
0|?
0L@
1&"
1T"
13#
03
1N
1d"
b0 T#
b0 $$
b0 R$
b0 "%
b0 P%
b0 ~%
b0 N&
b0 |&
b0 L'
b0 z'
b0 J(
b0 x(
b0 H)
b0 v)
b0 F*
b0 t*
b0 D+
b0 r+
b0 B,
b0 p,
b0 @-
b0 n-
b0 >.
b0 l.
b0 </
b0 j/
b0 :0
b0 h0
b0 81
b0 f1
b0 62
b0 d2
b0 43
b0 b3
b0 24
b0 `4
b0 05
b0 ^5
b0 .6
b0 \6
b0 ,7
b0 Z7
b0 *8
b0 X8
b0 (9
b0 V9
b0 &:
b0 T:
b0 $;
b0 R;
b0 "<
b0 P<
b0 ~<
b0 N=
b0 |=
b0 L>
b0 z>
b0 J?
b0 x?
b0 H@
b11 ""
1z"
0G#
b10 N#
0u#
b10 |#
0E$
b10 L$
0s$
b10 z$
0C%
b10 J%
0q%
b10 x%
0A&
b10 H&
0o&
b10 v&
0?'
b10 F'
0m'
b10 t'
0=(
b10 D(
0k(
b10 r(
0;)
b10 B)
0i)
b10 p)
09*
b10 @*
0g*
b10 n*
07+
b10 >+
0e+
b10 l+
05,
b10 <,
0c,
b10 j,
03-
b10 :-
0a-
b10 h-
01.
b10 8.
0_.
b10 f.
0//
b10 6/
0]/
b10 d/
0-0
b10 40
0[0
b10 b0
0+1
b10 21
0Y1
b10 `1
0)2
b10 02
0W2
b10 ^2
0'3
b10 .3
0U3
b10 \3
0%4
b10 ,4
0S4
b10 Z4
0#5
b10 *5
0Q5
b10 X5
0!6
b10 (6
0O6
b10 V6
0}6
b10 &7
0M7
b10 T7
0{7
b10 $8
0K8
b10 R8
0y8
b10 "9
0I9
b10 P9
0w9
b10 ~9
0G:
b10 N:
0u:
b10 |:
0E;
b10 L;
0s;
b10 z;
0C<
b10 J<
0q<
b10 x<
0A=
b10 H=
0o=
b10 v=
0?>
b10 F>
0m>
b10 t>
0=?
b10 D?
0k?
b10 r?
0;@
b10 B@
0B
0z
1{
1K"
1H#
b10 <#
b10 K#
1v#
b10 j#
b10 y#
1F$
b10 :$
b10 I$
1t$
b10 h$
b10 w$
1D%
b10 8%
b10 G%
1r%
b10 f%
b10 u%
1B&
b10 6&
b10 E&
1p&
b10 d&
b10 s&
1@'
b10 4'
b10 C'
1n'
b10 b'
b10 q'
1>(
b10 2(
b10 A(
1l(
b10 `(
b10 o(
1<)
b10 0)
b10 ?)
1j)
b10 ^)
b10 m)
1:*
b10 .*
b10 =*
1h*
b10 \*
b10 k*
18+
b10 ,+
b10 ;+
1f+
b10 Z+
b10 i+
16,
b10 *,
b10 9,
1d,
b10 X,
b10 g,
14-
b10 (-
b10 7-
1b-
b10 V-
b10 e-
12.
b10 &.
b10 5.
1`.
b10 T.
b10 c.
10/
b10 $/
b10 3/
1^/
b10 R/
b10 a/
1.0
b10 "0
b10 10
1\0
b10 P0
b10 _0
1,1
b10 ~0
b10 /1
1Z1
b10 N1
b10 ]1
1*2
b10 |1
b10 -2
1X2
b10 L2
b10 [2
1(3
b10 z2
b10 +3
1V3
b10 J3
b10 Y3
1&4
b10 x3
b10 )4
1T4
b10 H4
b10 W4
1$5
b10 v4
b10 '5
1R5
b10 F5
b10 U5
1"6
b10 t5
b10 %6
1P6
b10 D6
b10 S6
1~6
b10 r6
b10 #7
1N7
b10 B7
b10 Q7
1|7
b10 p7
b10 !8
1L8
b10 @8
b10 O8
1z8
b10 n8
b10 }8
1J9
b10 >9
b10 M9
1x9
b10 l9
b10 {9
1H:
b10 <:
b10 K:
1v:
b10 j:
b10 y:
1F;
b10 :;
b10 I;
1t;
b10 h;
b10 w;
1D<
b10 8<
b10 G<
1r<
b10 f<
b10 u<
1B=
b10 6=
b10 E=
1p=
b10 d=
b10 s=
1@>
b10 4>
b10 C>
1n>
b10 b>
b10 q>
1>?
b10 2?
b10 A?
1l?
b10 `?
b10 o?
1<@
b10 0@
b10 ?@
0I
1p
1@"
1n"
1>#
1l#
1<$
1j$
1:%
1h%
18&
1f&
16'
1d'
14(
1b(
12)
1`)
10*
1^*
1.+
1\+
1,,
1Z,
1*-
1X-
1(.
1V.
1&/
1T/
1$0
1R0
1"1
1P1
1~1
1N2
1|2
1L3
1z3
1J4
1x4
1H5
1v5
1F6
1t6
1D7
1r7
1B8
1p8
1@9
1n9
1>:
1l:
1<;
1j;
1:<
1h<
18=
1f=
16>
1d>
14?
1b?
12@
0H
0v
1x
0F"
1H"
0t"
1v"
0D#
1F#
0r#
1t#
0B$
1D$
0p$
1r$
0@%
1B%
0n%
1p%
0>&
1@&
0l&
1n&
0<'
1>'
0j'
1l'
0:(
1<(
0h(
1j(
08)
1:)
0f)
1h)
06*
18*
0d*
1f*
04+
16+
0b+
1d+
02,
14,
0`,
1b,
00-
12-
0^-
1`-
0..
10.
0\.
1^.
0,/
1./
0Z/
1\/
0*0
1,0
0X0
1Z0
0(1
1*1
0V1
1X1
0&2
1(2
0T2
1V2
0$3
1&3
0R3
1T3
0"4
1$4
0P4
1R4
0~4
1"5
0N5
1P5
0|5
1~5
0L6
1N6
0z6
1|6
0J7
1L7
0x7
1z7
0H8
1J8
0v8
1x8
0F9
1H9
0t9
1v9
0D:
1F:
0r:
1t:
0B;
1D;
0p;
1r;
0@<
1B<
0n<
1p<
0>=
1@=
0l=
1n=
0<>
1>>
0j>
1l>
0:?
1<?
0h?
1j?
08@
1:@
17
18
1d
14"
1b"
12#
1`#
10$
1^$
1.%
1\%
1,&
1Z&
1*'
1X'
1((
1V(
1&)
1T)
1$*
1R*
1"+
1P+
1~+
1N,
1|,
1L-
1z-
1J.
1x.
1H/
1v/
1F0
1t0
1D1
1r1
1B2
1p2
1@3
1n3
1>4
1l4
1<5
1j5
1:6
1h6
187
1f7
168
1d8
149
1b9
12:
1`:
10;
1^;
1.<
1\<
1,=
1Z=
1*>
1X>
1(?
1V?
1&@
b110 !
b110 *
b110 0
b110 /
0$
1i
12"
0;
1c"
19"
0g"
b110 #
b110 2
0b
1)"
b11 !"
b11 ."
16"
1`"
00#
1,"
0L"
0Y
15"
1W"
b11 O"
b11 \"
0'#
b0 }"
b0 ,#
0\
b1 ("
1f
0S
b0 Q
b0 ^
1Z"
0*#
1y
b111 n
b111 }
0|
0V
b0 X
1e
b1 V"
b0 &#
0K
19
b1111111111111111111111111111111111111111111111111111111111111111 1
b10 R
1I"
b11 P"
0w"
b10 ~"
1L
0M
b10 @
b10 O
0J"
b111 >"
b111 M"
1x"
b10 l"
b10 {"
1A
1?"
0m"
1E
1C"
0q"
b1 >
b1 C
1<
b1 <"
b1 A"
1:"
b10 j"
b10 o"
0h"
b101000 '
b101000 .
b10011111000101000 +
b111 (
b111 4
#30
